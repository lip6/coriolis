* Spice description of inv_x2
* Spice driver version 1363757992
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:43

* INTERF i nq vdd vss 


.subckt inv_x2 1 3 2 4 
* NET 1 = i
* NET 2 = vdd
* NET 3 = nq
* NET 4 = vss
Mtr_00002 3 1 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00001 4 1 3 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C4 1 4 8.60287e-16
C3 2 4 1.04191e-15
C2 3 4 1.22684e-15
C1 4 4 8.75833e-16
.ends inv_x2

