* Spice description of a2_x4
* Spice driver version 83533595
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:10

* INTERF i0 i1 q vdd vss 


.subckt a2_x4 4 3 2 1 7 
* NET 1 = vdd
* NET 2 = q
* NET 3 = i1
* NET 4 = i0
* NET 7 = vss
Xtr_00008 1 6 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 2 6 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 1 3 6 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00005 6 4 1 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00004 7 6 2 7 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 2 6 7 7 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 7 3 5 7 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 5 4 6 7 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C7 1 7 2.4749e-15
C6 2 7 1.08178e-15
C5 3 7 2.41961e-14
C4 4 7 1.8952e-14
C2 6 7 3.58946e-14
C1 7 7 1.83543e-15
.ends a2_x4

