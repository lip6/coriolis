* Spice description of buf_x8
* Spice driver version 2057223963
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:14

* INTERF i q vdd vss 


.subckt buf_x8 3 2 1 4 
* NET 1 = vdd
* NET 2 = q
* NET 3 = i
* NET 4 = vss
Xtr_00010 2 5 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 1 5 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 1 5 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 2 5 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 1 3 5 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00005 2 5 4 4 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 4 5 2 4 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 4 5 2 4 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 2 5 4 4 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 4 3 5 4 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C5 1 4 3.16371e-15
C4 2 4 3.29763e-15
C3 3 4 1.98449e-14
C2 4 4 2.38705e-15
C1 5 4 8.3284e-14
.ends buf_x8

