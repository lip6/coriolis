* Spice description of no2_x4
* Spice driver version 1024228264
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:58

* INTERF i0 i1 nq vdd vss 


.subckt no2_x4 1 2 7 5 8 
* NET 1 = i0
* NET 2 = i1
* NET 5 = vdd
* NET 7 = nq
* NET 8 = vss
Mtr_00010 5 6 3 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00009 7 3 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00008 5 3 7 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00007 5 2 4 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00006 4 1 6 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 3 6 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00004 8 3 7 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 7 3 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 6 2 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00001 8 1 6 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
C8 1 8 9.24715e-16
C7 2 8 8.17567e-16
C6 3 8 1.99373e-15
C4 5 8 2.51249e-15
C3 6 8 2.76016e-15
C2 7 8 1.22684e-15
C1 8 8 2.42677e-15
.ends no2_x4

