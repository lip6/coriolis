* Spice description of noa2ao222_x1
* Spice driver version -1590604005
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:24

* INTERF i0 i1 i2 i3 i4 nq vdd vss 


.subckt noa2ao222_x1 10 9 5 4 6 7 3 12 
* NET 3 = vdd
* NET 4 = i3
* NET 5 = i2
* NET 6 = i4
* NET 7 = nq
* NET 9 = i1
* NET 10 = i0
* NET 12 = vss
Xtr_00010 2 4 1 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 1 5 7 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 7 6 2 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 2 9 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 3 10 2 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00005 8 4 12 12 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Xtr_00004 12 5 8 12 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Xtr_00003 8 6 7 12 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Xtr_00002 7 9 11 12 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Xtr_00001 11 10 12 12 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
C11 2 12 9.70324e-16
C10 3 12 1.79971e-15
C9 4 12 1.6245e-14
C8 5 12 1.8135e-14
C7 6 12 1.69143e-14
C6 7 12 1.72074e-15
C5 8 12 4.45309e-16
C4 9 12 1.719e-14
C3 10 12 1.2224e-14
C1 12 12 2.1056e-15
.ends noa2ao222_x1

