* Spice description of nts_x2
* Spice driver version -335233253
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:26

* INTERF cmd i nq vdd vss 


.subckt nts_x2 5 8 6 3 10 
* NET 3 = vdd
* NET 5 = cmd
* NET 6 = nq
* NET 8 = i
* NET 10 = vss
Xtr_00010 3 8 1 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 4 5 3 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00008 2 8 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 6 4 2 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 1 4 6 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00005 4 5 10 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00004 10 8 7 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 9 8 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 6 5 9 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 7 5 6 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C8 3 10 2.44035e-15
C7 4 10 1.77683e-14
C6 5 10 3.37537e-14
C5 6 10 1.99345e-15
C3 8 10 4.38962e-14
C1 10 10 2.05203e-15
.ends nts_x2

