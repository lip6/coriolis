* Spice description of nxr2_x4
* Spice driver version -378462437
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:26

* INTERF i0 i1 nq vdd vss 


.subckt nxr2_x4 9 5 3 2 10 
* NET 2 = vdd
* NET 3 = nq
* NET 5 = i1
* NET 9 = i0
* NET 10 = vss
Xtr_00016 2 8 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00015 3 8 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00014 2 5 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 1 11 8 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 1 9 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 8 4 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 4 5 2 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00009 2 9 11 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00008 10 8 3 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00007 3 8 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00006 4 5 10 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00005 10 9 11 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00004 7 11 8 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 10 4 7 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 8 5 6 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 6 9 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C11 1 10 4.7288e-16
C10 2 10 4.06914e-15
C9 3 10 1.93831e-15
C8 4 10 2.84373e-14
C7 5 10 2.64414e-14
C4 8 10 4.33976e-14
C3 9 10 2.41345e-14
C2 10 10 3.30443e-15
C1 11 10 3.00018e-14
.ends nxr2_x4

