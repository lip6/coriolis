* Spice description of na2_x4
* Spice driver version 1444142875
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:17

* INTERF i0 i1 nq vdd vss 


.subckt na2_x4 6 5 3 1 4 
* NET 1 = vdd
* NET 3 = nq
* NET 4 = vss
* NET 5 = i1
* NET 6 = i0
Xtr_00010 1 5 8 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00009 8 6 1 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00008 3 2 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 1 2 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 2 8 1 1 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00005 4 5 7 4 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00004 7 6 8 4 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00003 3 2 4 4 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00002 2 8 4 4 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Xtr_00001 4 2 3 4 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
C8 1 4 2.06581e-15
C7 2 4 4.33156e-14
C6 3 4 1.66143e-15
C5 4 4 2.03707e-15
C4 5 4 1.8559e-14
C3 6 4 1.8559e-14
C1 8 4 1.79825e-14
.ends na2_x4

