* Spice description of xr2_x1
* Spice driver version 1355063067
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:34

* INTERF i0 i1 q vdd vss 


.subckt xr2_x1 8 4 7 2 10 
* NET 2 = vdd
* NET 4 = i1
* NET 7 = q
* NET 8 = i0
* NET 10 = vss
Xtr_00012 3 4 2 2 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00011 2 4 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 1 9 7 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 7 3 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 1 8 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 2 8 9 2 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00006 5 9 7 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 10 3 5 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 3 4 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 6 8 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 7 4 6 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 10 8 9 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C10 1 10 1.03148e-15
C9 2 10 2.08674e-15
C8 3 10 2.63298e-14
C7 4 10 3.49155e-14
C4 7 10 1.90461e-15
C3 8 10 2.7654e-14
C2 9 10 2.85741e-14
C1 10 10 2.08674e-15
.ends xr2_x1

