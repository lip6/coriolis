* Spice description of nts_x2
* Spice driver version 974969768
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:11

* INTERF cmd i nq vdd vss 


.subckt nts_x2 1 2 7 5 9 
* NET 1 = cmd
* NET 2 = i
* NET 5 = vdd
* NET 7 = nq
* NET 9 = vss
Mtr_00010 8 1 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00009 3 2 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.34U AS=0.6786P AD=0.6786P PS=5.26U PD=5.26U 
Mtr_00008 7 8 3 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.34U AS=0.6786P AD=0.6786P PS=5.26U PD=5.26U 
Mtr_00007 4 8 7 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.34U AS=0.6786P AD=0.6786P PS=5.26U PD=5.26U 
Mtr_00006 5 2 4 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.34U AS=0.6786P AD=0.6786P PS=5.26U PD=5.26U 
Mtr_00005 6 2 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.14U AS=0.3306P AD=0.3306P PS=2.86U PD=2.86U 
Mtr_00004 7 1 6 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.14U AS=0.3306P AD=0.3306P PS=2.86U PD=2.86U 
Mtr_00003 9 1 8 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00002 10 2 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.14U AS=0.3306P AD=0.3306P PS=2.86U PD=2.86U 
Mtr_00001 7 1 10 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.14U AS=0.3306P AD=0.3306P PS=2.86U PD=2.86U 
C10 1 9 1.55285e-15
C9 2 9 1.54897e-15
C6 5 9 2.41767e-15
C4 7 9 1.70901e-15
C3 8 9 2.21365e-15
C2 9 9 1.96765e-15
.ends nts_x2

