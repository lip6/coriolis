* Spice description of o4_x4
* Spice driver version 1147682587
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:28

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt o4_x4 7 10 8 6 5 1 11 
* NET 1 = vdd
* NET 5 = q
* NET 6 = i3
* NET 7 = i0
* NET 8 = i2
* NET 10 = i1
* NET 11 = vss
Xtr_00012 5 9 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 1 9 5 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 1 6 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 2 8 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 4 7 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 3 10 9 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 5 9 11 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 11 9 5 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 11 6 9 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 9 8 11 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 11 7 9 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 9 10 11 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C11 1 11 2.51826e-15
C7 5 11 2.04386e-15
C6 6 11 1.53915e-14
C5 7 11 1.53152e-14
C4 8 11 1.63711e-14
C3 9 11 2.30545e-14
C2 10 11 1.53152e-14
C1 11 11 2.19936e-15
.ends o4_x4

