* Spice description of sff1r_x4
* Spice driver version -1876422885
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:33

* INTERF ck i nrst q vdd vss 


.subckt sff1r_x4 17 14 7 5 4 18 
* NET 4 = vdd
* NET 5 = q
* NET 7 = nrst
* NET 9 = sff_s
* NET 10 = y
* NET 11 = sff_m
* NET 14 = i
* NET 15 = ckr
* NET 17 = ck
* NET 18 = vss
* NET 19 = nckr
Xtr_00028 5 9 4 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00027 9 15 1 4 sg13_lv_pmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Xtr_00026 4 9 5 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00025 1 5 4 4 sg13_lv_pmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Xtr_00024 10 19 9 4 sg13_lv_pmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Xtr_00023 4 7 10 4 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00022 11 19 3 4 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00021 3 10 4 4 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00020 10 11 4 4 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00019 2 15 11 4 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00018 4 16 2 4 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00017 16 14 4 4 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00016 4 19 15 4 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00015 19 17 4 4 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00014 13 15 11 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00013 11 19 12 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00012 18 9 5 18 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00011 5 9 18 18 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00010 18 5 6 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00009 6 19 9 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00008 9 15 10 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00007 10 7 8 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00006 8 11 18 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00005 18 10 13 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00004 12 16 18 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00003 18 17 19 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 15 19 18 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 18 14 16 18 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C16 4 18 5.21376e-15
C15 5 18 2.123e-14
C13 7 18 2.20053e-14
C11 9 18 3.47422e-14
C10 10 18 2.30769e-14
C9 11 18 3.6015e-14
C6 14 18 1.59913e-14
C5 15 18 7.76489e-14
C4 16 18 2.74223e-14
C3 17 18 1.9047e-14
C2 18 18 4.83623e-15
C1 19 18 1.01179e-13
.ends sff1r_x4

