* Spice description of no4_x1
* Spice driver version -7042136
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:01

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt no4_x1 4 1 3 2 9 7 10 
* NET 1 = i1
* NET 2 = i3
* NET 3 = i2
* NET 4 = i0
* NET 7 = vdd
* NET 9 = nq
* NET 10 = vss
Mtr_00008 8 4 9 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00007 7 2 5 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00006 5 3 6 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 6 1 8 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00004 9 1 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00003 9 2 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00002 10 3 9 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00001 10 4 9 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
C10 1 10 9.24715e-16
C9 2 10 9.24715e-16
C8 3 10 9.24715e-16
C7 4 10 8.17567e-16
C4 7 10 1.55138e-15
C2 9 10 2.26082e-15
C1 10 10 1.87818e-15
.ends no4_x1

