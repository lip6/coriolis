* Spice description of mx2_x4
* Spice driver version -375185637
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:15

* INTERF cmd i0 i1 q vdd vss 


.subckt mx2_x4 9 10 5 4 3 11 
* NET 3 = vdd
* NET 4 = q
* NET 5 = i1
* NET 9 = cmd
* NET 10 = i0
* NET 11 = vss
Xtr_00014 4 7 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 3 5 2 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00012 1 10 3 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00011 3 9 12 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00010 2 12 7 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00009 7 9 1 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00008 3 7 4 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 11 5 6 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00006 6 9 7 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00005 7 12 8 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00004 8 10 11 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00003 11 9 12 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 4 7 11 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 11 7 4 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C10 3 11 3.87147e-15
C9 4 11 1.93831e-15
C8 5 11 2.12638e-14
C6 7 11 4.32593e-14
C4 9 11 5.39741e-14
C3 10 11 1.7193e-14
C2 11 11 3.02522e-15
C1 12 11 1.60395e-14
.ends mx2_x4

