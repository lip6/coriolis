* Spice description of on12_x4
* Spice driver version -1533351000
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:27

* INTERF i0 i1 q vdd vss 


.subckt on12_x4 1 4 7 5 8 
* NET 1 = i0
* NET 4 = i1
* NET 5 = vdd
* NET 7 = q
* NET 8 = vss
Mtr_00010 2 3 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00009 6 4 2 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00008 5 1 3 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.02U AS=0.2958P AD=0.2958P PS=2.62U PD=2.62U 
Mtr_00007 5 6 7 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00006 7 6 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 6 4 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00004 8 3 6 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00003 3 1 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.54U AS=0.1566P AD=0.1566P PS=1.66U PD=1.66U 
Mtr_00002 8 6 7 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 7 6 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C8 1 8 1.27591e-15
C6 3 8 1.6097e-15
C5 4 8 1.57438e-15
C4 5 8 3.44842e-15
C3 6 8 2.43977e-15
C2 7 8 1.22684e-15
C1 8 8 3.05197e-15
.ends on12_x4

