* Spice description of na4_x4
* Spice driver version 1928847131
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:18

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt na4_x4 5 6 3 2 9 1 11 
* NET 1 = vdd
* NET 2 = i3
* NET 3 = i2
* NET 5 = i0
* NET 6 = i1
* NET 9 = nq
* NET 11 = vss
Xtr_00014 1 12 9 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 9 12 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 1 10 12 1 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00011 10 5 1 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00010 1 6 10 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00009 10 3 1 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00008 1 2 10 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00007 11 12 9 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00006 9 12 11 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 11 10 12 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 8 5 11 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 7 6 8 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 10 2 4 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 4 3 7 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C12 1 11 2.43007e-15
C11 2 11 1.95386e-14
C10 3 11 2.09464e-14
C8 5 11 1.95386e-14
C7 6 11 1.98905e-14
C4 9 11 2.05734e-15
C3 10 11 1.52642e-14
C2 11 11 2.31745e-15
C1 12 11 4.72809e-14
.ends na4_x4

