* Spice description of inv_x1
* Spice driver version 212172571
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:14

* INTERF i nq vdd vss 


.subckt inv_x1 2 4 1 3 
* NET 1 = vdd
* NET 2 = i
* NET 3 = vss
* NET 4 = nq
Xtr_00002 4 2 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00001 4 2 3 3 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C4 1 3 1.08664e-15
C3 2 3 2.00735e-14
C2 3 3 1.07285e-15
C1 4 3 1.93831e-15
.ends inv_x1

