* Spice description of oa3ao322_x2
* Spice driver version 264706984
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:25

* INTERF i0 i1 i2 i3 i4 i5 i6 q vdd vss 


.subckt oa3ao322_x2 11 10 9 1 4 3 2 16 12 17 
* NET 1 = i3
* NET 2 = i6
* NET 3 = i5
* NET 4 = i4
* NET 9 = i2
* NET 10 = i1
* NET 11 = i0
* NET 12 = vdd
* NET 16 = q
* NET 17 = vss
Mtr_00016 16 15 12 12 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00015 5 3 7 12 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00014 5 4 6 12 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00013 12 11 7 12 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.435P AD=0.435P PS=3.58U PD=3.58U 
Mtr_00012 7 10 12 12 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.435P AD=0.435P PS=3.58U PD=3.58U 
Mtr_00011 12 9 7 12 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.435P AD=0.435P PS=3.58U PD=3.58U 
Mtr_00010 7 2 15 12 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.435P AD=0.435P PS=3.58U PD=3.58U 
Mtr_00009 6 1 15 12 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00008 17 15 16 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00007 15 9 13 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.14U AS=0.3306P AD=0.3306P PS=2.86U PD=2.86U 
Mtr_00006 8 4 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.54U AS=0.1566P AD=0.1566P PS=1.66U PD=1.66U 
Mtr_00005 13 10 14 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.14U AS=0.3306P AD=0.3306P PS=2.86U PD=2.86U 
Mtr_00004 14 11 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.14U AS=0.3306P AD=0.3306P PS=2.86U PD=2.86U 
Mtr_00003 17 1 8 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.54U AS=0.1566P AD=0.1566P PS=1.66U PD=1.66U 
Mtr_00002 8 2 15 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.54U AS=0.1566P AD=0.1566P PS=1.66U PD=1.66U 
Mtr_00001 17 3 8 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.54U AS=0.1566P AD=0.1566P PS=1.66U PD=1.66U 
C17 1 17 9.66594e-16
C16 2 17 7.48234e-16
C15 3 17 1.04475e-15
C14 4 17 9.39915e-16
C11 7 17 1.49471e-15
C10 8 17 9.42902e-16
C9 9 17 1.07273e-15
C8 10 17 9.76258e-16
C7 11 17 8.42431e-16
C6 12 17 2.64694e-15
C3 15 17 2.78895e-15
C2 16 17 1.22684e-15
C1 17 17 2.7273e-15
.ends oa3ao322_x2

