* Spice description of zero_x0
* Spice driver version -381326424
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:33

* INTERF nq vdd vss 


.subckt zero_x0 2 1 3 
* NET 1 = vdd
* NET 2 = nq
* NET 3 = vss
Mtr_00001 2 1 3 3 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.1218P AD=0.1218P PS=1.42U PD=1.42U 
C3 1 3 1.76813e-15
C2 2 3 9.32188e-16
C1 3 3 8.75833e-16
.ends zero_x0

