* Spice description of noa2a2a2a24_x4
* Spice driver version -108110053
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:24

* INTERF i0 i1 i2 i3 i4 i5 i6 i7 nq vdd vss 


.subckt noa2a2a2a24_x4 6 7 10 11 13 14 17 18 9 2 20 
* NET 2 = vdd
* NET 6 = i0
* NET 7 = i1
* NET 9 = nq
* NET 10 = i2
* NET 11 = i3
* NET 13 = i4
* NET 14 = i5
* NET 17 = i6
* NET 18 = i7
* NET 20 = vss
Xtr_00022 5 15 2 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00021 2 5 9 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00020 9 5 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00019 2 6 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00018 1 7 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00017 3 10 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00016 1 11 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00015 3 13 4 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00014 4 14 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 4 17 15 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 15 18 4 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 5 15 20 20 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00010 20 5 9 20 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00009 9 5 20 20 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00008 20 6 8 20 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00007 8 7 15 20 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00006 20 10 12 20 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 12 11 15 20 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 15 13 16 20 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 16 14 20 20 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 15 17 19 20 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 19 18 20 20 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C20 1 20 7.52081e-16
C19 2 20 4.51629e-15
C18 3 20 9.61383e-16
C17 4 20 9.61383e-16
C16 5 20 2.9742e-14
C15 6 20 1.47638e-14
C14 7 20 1.54677e-14
C12 9 20 2.48991e-15
C11 10 20 1.47638e-14
C10 11 20 1.51158e-14
C8 13 20 1.47638e-14
C7 14 20 1.47638e-14
C6 15 20 2.02278e-14
C4 17 20 1.47638e-14
C3 18 20 1.50395e-14
C1 20 20 3.63995e-15
.ends noa2a2a2a24_x4

