* Spice description of nao2o22_x1
* Spice driver version 990751656
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:53

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt nao2o22_x1 4 3 2 1 8 7 10 
* NET 1 = i3
* NET 2 = i2
* NET 3 = i1
* NET 4 = i0
* NET 7 = vdd
* NET 8 = nq
* NET 10 = vss
Mtr_00008 6 1 8 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00007 7 2 6 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00006 8 3 5 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 5 4 7 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00004 10 2 9 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 9 1 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 8 3 9 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 9 4 8 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C10 1 10 9.67435e-16
C9 2 10 8.038e-16
C8 3 10 8.60287e-16
C7 4 10 9.92572e-16
C4 7 10 1.63174e-15
C3 8 10 1.30721e-15
C2 9 10 1.25899e-15
C1 10 10 1.3853e-15
.ends nao2o22_x1

