* Spice description of buf_x4
* Spice driver version -213722200
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:40

* INTERF i q vdd vss 


.subckt buf_x4 1 4 2 5 
* NET 1 = i
* NET 2 = vdd
* NET 4 = q
* NET 5 = vss
Mtr_00006 2 3 4 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 2 1 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00004 4 3 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00003 4 3 5 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 3 1 5 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00001 5 3 4 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C5 1 5 9.7156e-16
C4 2 5 2.00302e-15
C3 3 5 2.34697e-15
C2 4 5 1.22684e-15
C1 5 5 1.67086e-15
.ends buf_x4

