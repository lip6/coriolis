* Spice description of a3_x4
* Spice driver version 2105387944
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:33

* INTERF i0 i1 i2 q vdd vss 


.subckt a3_x4 4 2 1 9 5 8 
* NET 1 = i2
* NET 2 = i1
* NET 4 = i0
* NET 5 = vdd
* NET 8 = vss
* NET 9 = q
Mtr_00010 5 2 3 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00009 3 1 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00008 3 4 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00007 5 3 9 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00006 9 3 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 9 3 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00004 6 1 3 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 7 2 6 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 8 4 7 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 8 3 9 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C9 1 8 1.06324e-15
C8 2 8 1.01428e-15
C7 3 8 3.07916e-15
C6 4 8 7.39551e-16
C5 5 8 2.47124e-15
C2 8 8 2.01051e-15
C1 9 8 1.93938e-15
.ends a3_x4

