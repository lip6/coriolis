* Spice description of noa2a22_x4
* Spice driver version -1866387685
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:23

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt noa2a22_x4 10 9 6 5 3 2 12 
* NET 2 = vdd
* NET 3 = nq
* NET 5 = i3
* NET 6 = i2
* NET 9 = i1
* NET 10 = i0
* NET 12 = vss
Xtr_00014 1 9 7 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00013 7 10 1 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00012 3 4 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 2 4 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 2 7 4 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00009 1 6 2 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00008 2 5 1 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00007 7 9 11 12 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00006 11 10 12 12 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00005 3 4 12 12 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 12 4 3 12 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 12 7 4 12 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 8 5 7 12 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 12 6 8 12 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C12 1 12 8.6004e-16
C11 2 12 3.78095e-15
C10 3 12 1.99345e-15
C9 4 12 3.13076e-14
C8 5 12 2.4894e-14
C7 6 12 2.13745e-14
C6 7 12 2.15407e-14
C4 9 12 1.8559e-14
C3 10 12 1.83108e-14
C1 12 12 3.58223e-15
.ends noa2a22_x4

