* Spice description of o2_x2
* Spice driver version 597941160
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:13

* INTERF i0 i1 q vdd vss 


.subckt o2_x2 1 2 6 4 7 
* NET 1 = i0
* NET 2 = i1
* NET 4 = vdd
* NET 6 = q
* NET 7 = vss
Mtr_00006 4 1 3 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 3 2 5 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00004 6 5 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00003 7 2 5 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00002 5 1 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00001 6 5 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C7 1 7 7.3965e-16
C6 2 7 1.01861e-15
C4 4 7 1.21548e-15
C3 5 7 2.17821e-15
C2 6 7 1.22684e-15
C1 7 7 1.52085e-15
.ends o2_x2

