CARACTERISATION_OTA_CASCODE_SIMPLE_REPLIE

* alimentations *
vdd evdd 0 3.300000
vss evss 0 0.000000
gfoncd evdd 0 evdd 0 1.0e-15

* acces aux modeles de simulation *
.include /users/cao/porte/OCEAN/oceane/share/envtech/modeles/proprietaires/ams0.35/eldo_bsim3v3 

* dispositif principal *

.SUBCKT OTACSRND1 ep em sp evp1 evp2 evc1 evc3 evdd evss
*infoceane:netpolar evp1 evp2 evc1 evc3
MN1 nbi1c_1 ep 2_1 evss modn_typ W=1.75000u L=1.95000u M=10
+ ad=1.066p as=2.132p pd=2.977u ps=5.954u
+ nrs=0.000 nrd=0.000 
MN2 nbi2c_1 em 2_1 evss modn_typ W=1.75000u L=1.95000u M=10
+ ad=1.066p as=2.132p pd=2.977u ps=5.954u
+ nrs=0.000 nrd=0.000 
MN5 2_1 evp1 evss evss modn_typ W=4.45000u L=2.65000u M=12
+ ad=2.686p as=5.372p pd=5.677u ps=11.354u
+ nrs=0.000 nrd=0.000 
MP1C ndm1c_1 evc1 nbi1c_1 nbi1c_1 modp_typ W=8.45000u L=1.95000u M=6
+ ad=5.093p as=10.186p pd=9.688u ps=19.377u
+ nrs=0.000 nrd=0.000 
D_MP1C evss nbi1c_1 dwell_sub AREA=113.295p PJ=43.100u 
MP2C sp evc1 nbi2c_1 nbi2c_1 modp_typ W=8.45000u L=1.95000u M=6
+ ad=5.093p as=10.186p pd=9.688u ps=19.377u
+ nrs=0.000 nrd=0.000 
D_MP2C evss nbi2c_1 dwell_sub AREA=113.295p PJ=43.100u 
MP7 nbi1c_1 evp2 evdd evdd modp_typ W=17.40000u L=1.95000u M=6
+ ad=10.463p as=20.926p pd=18.638u ps=37.277u
+ nrs=0.000 nrd=0.000 
D_MP7 evss evdd dwell_sub AREA=194.740p PJ=61.000u 
MP8 nbi2c_1 evp2 evdd evdd modp_typ W=17.40000u L=1.95000u M=6
+ ad=10.463p as=20.926p pd=18.638u ps=37.277u
+ nrs=0.000 nrd=0.000 
D_MP8 evss evdd dwell_sub AREA=194.740p PJ=61.000u 
MN3 nbi3c_1 ndm1c_1 evss evss modn_typ W=0.50000u L=2.65000u M=2
+ ad=0.316p as=0.474p pd=1.727u ps=2.590u
+ nrs=0.000 nrd=0.000 
MN4 nbi4c_1 ndm1c_1 evss evss modn_typ W=0.50000u L=2.65000u M=2
+ ad=0.316p as=0.474p pd=1.727u ps=2.590u
+ nrs=0.000 nrd=0.000 
MN3C ndm1c_1 evc3 nbi3c_1 evss modn_typ W=1.75000u L=1.95000u M=10
+ ad=1.066p as=2.132p pd=2.977u ps=5.954u
+ nrs=0.000 nrd=0.000 
MN4C sp evc3 nbi4c_1 evss modn_typ W=1.75000u L=1.95000u M=10
+ ad=1.066p as=2.132p pd=2.977u ps=5.954u
+ nrs=0.000 nrd=0.000 
.ENDS OTACSRND1
*
XOTACSRND1 ep em sp evp1 evp2 evc1 evc3 evdd evss OTACSRND1
*

* dispositif auxiliaire 1 *
.SUBCKT POLAR_OTACSRND1 evp1 evp2 evc1 evc3 evdd evss
vp1 evp1 0 0.6830
vp2 evp2 0 2.4598
vc1 evc1 0 2.1580
vc3 evc3 0 1.8255
rfonc_vdd evdd 0 1.0e15 
rfonc_vss evss 0 1.0e15 
.ENDS POLAR_OTACSRND1
*
XPOLAR_OTACSRND1 evp1 evp2 evc1 evc3 evdd evss POLAR_OTACSRND1
*

* dispositif auxiliaire 3 *
.SUBCKT CHARGE_OTACSRND1 sp smc
CL sp smc 3.000000e-12
.ENDS CHARGE_OTACSRND1
*
XCHARGE_OTACSRND1 sp smc CHARGE_OTACSRND1
*

* mode commun en entree *
vemc emc 0 1.650000

* mode commun en sortie *
vsmc smc 0 1.650000

* determination des points de repos *
vcct sp em dc 0.000000
vop ep emc dc 0.0
.op

* options de simulation *
.option nowavecomplex stat=3 nomod analog eps=1.0e-6 numdgt=8

* temperature de simulation *
.temp 27.00

.nodeset v(sp)=1.650000


* fin de fichier *
.end

