* Spice description of nao22_x4
* Spice driver version -333807845
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:18

* INTERF i0 i1 i2 nq vdd vss 


.subckt nao22_x4 6 5 8 4 2 10 
* NET 2 = vdd
* NET 4 = nq
* NET 5 = i1
* NET 6 = i0
* NET 8 = i2
* NET 10 = vss
Xtr_00012 2 3 4 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 4 3 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 1 5 7 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00009 2 6 1 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00008 7 8 2 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00007 2 7 3 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00006 4 3 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 10 3 4 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 7 5 9 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00003 9 8 10 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 9 6 7 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 10 7 3 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C9 2 10 3.87331e-15
C8 3 10 4.01623e-14
C7 4 10 1.99345e-15
C6 5 10 2.70914e-14
C5 6 10 2.60261e-14
C4 7 10 1.64383e-14
C3 8 10 2.27061e-14
C2 9 10 5.00451e-16
C1 10 10 3.03967e-15
.ends nao22_x4

