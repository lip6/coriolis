* Spice description of oa22_x4
* Spice driver version 709237672
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:18

* INTERF i0 i1 i2 q vdd vss 


.subckt oa22_x4 2 4 3 6 5 9 
* NET 2 = i0
* NET 3 = i2
* NET 4 = i1
* NET 5 = vdd
* NET 6 = q
* NET 9 = vss
Mtr_00010 5 8 6 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00009 6 8 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00008 1 4 8 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00007 5 3 1 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00006 8 2 1 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00005 6 8 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00004 6 8 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 9 2 7 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00002 7 4 8 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00001 8 3 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
C9 1 9 6.5896e-16
C8 2 9 1.06968e-15
C7 3 9 9.61108e-16
C6 4 9 1.23481e-15
C5 5 9 3.05359e-15
C4 6 9 1.22684e-15
C2 8 9 2.15615e-15
C1 9 9 2.63571e-15
.ends oa22_x4

