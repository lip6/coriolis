* Spice description of na4_x1
* Spice driver version 62734107
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:17

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt na4_x1 8 7 2 3 6 1 10 
* NET 1 = vdd
* NET 2 = i2
* NET 3 = i3
* NET 6 = nq
* NET 7 = i1
* NET 8 = i0
* NET 10 = vss
Xtr_00008 1 3 6 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00007 1 7 6 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00006 6 8 1 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00005 6 2 1 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00004 6 3 4 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 4 2 5 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 9 8 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 5 7 9 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C10 1 10 1.87762e-15
C9 2 10 1.88347e-14
C8 3 10 1.96148e-14
C5 6 10 2.53966e-15
C4 7 10 1.88347e-14
C3 8 10 1.91866e-14
C1 10 10 1.569e-15
.ends na4_x1

