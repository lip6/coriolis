* Spice description of noa3ao322_x1
* Spice driver version -600080613
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:25

* INTERF i0 i1 i2 i3 i4 i5 i6 nq vdd vss 


.subckt noa3ao322_x1 14 13 9 5 6 7 8 10 4 16 
* NET 4 = vdd
* NET 5 = i3
* NET 6 = i4
* NET 7 = i5
* NET 8 = i6
* NET 9 = i2
* NET 10 = nq
* NET 13 = i1
* NET 14 = i0
* NET 16 = vss
Xtr_00014 10 8 3 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 3 9 4 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 4 13 3 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 3 14 4 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 2 5 10 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 1 6 2 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 3 7 1 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 11 8 10 16 sg13_lv_nmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
Xtr_00006 10 9 12 16 sg13_lv_nmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
Xtr_00005 12 13 15 16 sg13_lv_nmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
Xtr_00004 15 14 16 16 sg13_lv_nmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
Xtr_00003 16 5 11 16 sg13_lv_nmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
Xtr_00002 11 6 16 16 sg13_lv_nmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
Xtr_00001 16 7 11 16 sg13_lv_nmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
C14 3 16 1.17711e-15
C13 4 16 2.45714e-15
C12 5 16 1.1872e-14
C11 6 16 1.1872e-14
C10 7 16 1.1872e-14
C9 8 16 1.09687e-14
C8 9 16 1.1872e-14
C7 10 16 1.74831e-15
C6 11 16 4.86665e-16
C4 13 16 1.21477e-14
C3 14 16 1.15201e-14
C1 16 16 2.6875e-15
.ends noa3ao322_x1

