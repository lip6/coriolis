* Spice description of nxr2_x1
* Spice driver version 1740159912
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:12

* INTERF i0 i1 nq vdd vss 


.subckt nxr2_x1 3 1 8 4 7 
* NET 1 = i1
* NET 3 = i0
* NET 4 = vdd
* NET 7 = vss
* NET 8 = nq
Mtr_00012 4 2 5 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.34U AS=0.6786P AD=0.6786P PS=5.26U PD=5.26U 
Mtr_00011 5 6 8 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.34U AS=0.6786P AD=0.6786P PS=5.26U PD=5.26U 
Mtr_00010 8 1 5 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.34U AS=0.6786P AD=0.6786P PS=5.26U PD=5.26U 
Mtr_00009 5 3 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.34U AS=0.6786P AD=0.6786P PS=5.26U PD=5.26U 
Mtr_00008 2 1 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00007 4 3 6 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00006 10 1 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.14U AS=0.3306P AD=0.3306P PS=2.86U PD=2.86U 
Mtr_00005 8 6 10 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.14U AS=0.3306P AD=0.3306P PS=2.86U PD=2.86U 
Mtr_00004 9 2 8 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.14U AS=0.3306P AD=0.3306P PS=2.86U PD=2.86U 
Mtr_00003 7 3 9 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.14U AS=0.3306P AD=0.3306P PS=2.86U PD=2.86U 
Mtr_00002 6 3 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00001 7 1 2 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
C10 1 7 1.92291e-15
C9 2 7 2.18588e-15
C8 3 7 1.31112e-15
C7 4 7 2.14121e-15
C6 5 7 1.1947e-15
C5 6 7 1.57758e-15
C4 7 7 2.14121e-15
C3 8 7 1.78937e-15
.ends nxr2_x1

