* Spice description of na3_x1
* Spice driver version -1981023320
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:49

* INTERF i0 i1 i2 nq vdd vss 


.subckt na3_x1 2 3 4 6 1 5 
* NET 1 = vdd
* NET 2 = i0
* NET 3 = i1
* NET 4 = i2
* NET 5 = vss
* NET 6 = nq
Mtr_00006 6 4 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00005 1 3 6 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00004 6 2 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 7 4 6 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.62U AS=0.4698P AD=0.4698P PS=3.82U PD=3.82U 
Mtr_00002 5 2 8 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.62U AS=0.4698P AD=0.4698P PS=3.82U PD=3.82U 
Mtr_00001 8 3 7 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.62U AS=0.4698P AD=0.4698P PS=3.82U PD=3.82U 
C8 1 5 1.46192e-15
C7 2 5 1.05763e-15
C6 3 5 9.50487e-16
C5 4 5 9.50487e-16
C4 5 5 1.21548e-15
C3 6 5 1.96617e-15
.ends na3_x1

