* Spice description of ao2o22_x2
* Spice driver version -1532334309
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:13

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt ao2o22_x2 9 5 7 6 4 3 8 
* NET 3 = vdd
* NET 4 = q
* NET 5 = i1
* NET 6 = i3
* NET 7 = i2
* NET 8 = vss
* NET 9 = i0
Xtr_00010 3 6 1 3 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00009 10 5 2 3 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00008 4 10 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 1 7 10 3 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00006 2 9 3 3 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00005 10 9 11 8 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Xtr_00004 11 5 10 8 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Xtr_00003 4 10 8 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 11 6 8 8 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Xtr_00001 8 7 11 8 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
C9 3 8 2.46702e-15
C8 4 8 1.93831e-15
C7 5 8 1.81795e-14
C6 6 8 1.88558e-14
C5 7 8 2.37925e-14
C4 8 8 2.3241e-15
C3 9 8 1.79313e-14
C2 10 8 1.61079e-14
C1 11 8 8.18684e-16
.ends ao2o22_x2

