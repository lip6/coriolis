* Spice description of o3_x4
* Spice driver version -424849637
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:27

* INTERF i0 i1 i2 q vdd vss 


.subckt o3_x4 4 6 7 5 1 8 
* NET 1 = vdd
* NET 4 = i0
* NET 5 = q
* NET 6 = i1
* NET 7 = i2
* NET 8 = vss
Xtr_00010 1 4 2 1 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00009 2 6 3 1 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00008 3 7 9 1 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00007 1 9 5 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 5 9 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00005 8 4 9 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 9 6 8 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 8 7 9 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 8 9 5 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 5 9 8 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C9 1 8 2.4955e-15
C6 4 8 1.53915e-14
C5 5 8 1.99345e-15
C4 6 8 1.57434e-14
C3 7 8 1.50395e-14
C2 8 8 2.16348e-15
C1 9 8 4.0414e-14
.ends o3_x4

