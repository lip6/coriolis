* Spice description of no4_x4
* Spice driver version -229077221
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:22

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt no4_x4 7 10 8 9 6 1 12 
* NET 1 = vdd
* NET 6 = nq
* NET 7 = i0
* NET 8 = i2
* NET 9 = i3
* NET 10 = i1
* NET 12 = vss
Xtr_00014 2 7 3 1 sg13_lv_pmos L=0.13U W=3.02U AS=0.7248P AD=0.7248P PS=6.52U PD=6.52U 
Xtr_00013 4 8 2 1 sg13_lv_pmos L=0.13U W=3.02U AS=0.7248P AD=0.7248P PS=6.52U PD=6.52U 
Xtr_00012 1 9 4 1 sg13_lv_pmos L=0.13U W=3.02U AS=0.7248P AD=0.7248P PS=6.52U PD=6.52U 
Xtr_00011 5 11 1 1 sg13_lv_pmos L=0.13U W=1.59U AS=0.3816P AD=0.3816P PS=3.67U PD=3.67U 
Xtr_00010 1 5 6 1 sg13_lv_pmos L=0.13U W=3.02U AS=0.7248P AD=0.7248P PS=6.52U PD=6.52U 
Xtr_00009 6 5 1 1 sg13_lv_pmos L=0.13U W=3.02U AS=0.7248P AD=0.7248P PS=6.52U PD=6.52U 
Xtr_00008 3 10 11 1 sg13_lv_pmos L=0.13U W=3.02U AS=0.7248P AD=0.7248P PS=6.52U PD=6.52U 
Xtr_00007 12 5 6 12 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00006 6 5 12 12 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 11 10 12 12 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00004 11 8 12 12 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00003 12 9 11 12 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 12 7 11 12 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 5 11 12 12 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C12 1 12 3.30366e-15
C8 5 12 5.13782e-14
C7 6 12 1.74532e-15
C6 7 12 1.74269e-14
C5 8 12 1.60191e-14
C4 9 12 1.53152e-14
C3 10 12 1.63711e-14
C2 11 12 1.96921e-14
C1 12 12 2.64543e-15
.ends no4_x4

