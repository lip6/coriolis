* Spice description of oa2a2a23_x4
* Spice driver version -94044389
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:30

* INTERF i0 i1 i2 i3 i4 i5 q vdd vss 


.subckt oa2a2a23_x4 6 5 8 9 10 13 4 1 15 
* NET 1 = vdd
* NET 4 = q
* NET 5 = i1
* NET 6 = i0
* NET 8 = i2
* NET 9 = i3
* NET 10 = i4
* NET 13 = i5
* NET 15 = vss
Xtr_00016 1 12 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00015 4 12 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00014 1 6 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 2 5 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 12 13 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 3 8 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 2 9 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 3 10 12 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 15 12 4 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00007 4 12 15 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00006 7 5 12 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 15 8 11 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 14 13 15 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 15 6 7 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 11 9 12 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 12 10 14 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C15 1 15 4.05966e-15
C14 2 15 7.91783e-16
C13 3 15 7.49757e-16
C12 4 15 1.99345e-15
C11 5 15 2.04337e-14
C10 6 15 2.11376e-14
C8 8 15 2.04337e-14
C7 9 15 2.04337e-14
C6 10 15 1.9177e-14
C4 12 15 3.59026e-14
C3 13 15 2.04337e-14
C1 15 15 3.19779e-15
.ends oa2a2a23_x4

