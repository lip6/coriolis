* Spice description of noa2a2a23_x1
* Spice driver version -647590117
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:23

* INTERF i0 i1 i2 i3 i4 i5 nq vdd vss 


.subckt noa2a2a23_x1 5 4 8 7 11 12 10 1 14 
* NET 1 = vdd
* NET 4 = i1
* NET 5 = i0
* NET 7 = i3
* NET 8 = i2
* NET 10 = nq
* NET 11 = i4
* NET 12 = i5
* NET 14 = vss
Xtr_00012 10 12 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 3 11 10 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 2 7 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 3 8 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 1 5 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 2 4 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 9 7 10 14 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 14 8 9 14 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 6 4 10 14 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 14 5 6 14 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 10 11 13 14 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 13 12 14 14 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C14 1 14 2.72688e-15
C13 2 14 7.65866e-16
C12 3 14 7.49757e-16
C11 4 14 1.47638e-14
C10 5 14 1.47638e-14
C8 7 14 2.37121e-14
C7 8 14 2.25066e-14
C5 10 14 2.47172e-15
C4 11 14 2.51924e-14
C3 12 14 1.86241e-14
C1 14 14 2.42542e-15
.ends noa2a2a23_x1

