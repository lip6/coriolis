* Spice description of noa2a2a23_x4
* Spice driver version 1658261275
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:23

* INTERF i0 i1 i2 i3 i4 i5 nq vdd vss 


.subckt noa2a2a23_x4 6 7 11 10 9 15 5 1 16 
* NET 1 = vdd
* NET 5 = nq
* NET 6 = i0
* NET 7 = i1
* NET 9 = i4
* NET 10 = i3
* NET 11 = i2
* NET 15 = i5
* NET 16 = vss
Xtr_00018 1 6 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00017 14 15 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00016 3 9 14 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00015 2 10 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00014 3 11 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 1 4 5 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 5 4 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 2 7 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 4 14 1 1 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00009 16 6 8 16 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00008 13 15 16 16 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00007 14 9 13 16 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00006 12 10 14 16 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 16 11 12 16 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 16 4 5 16 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 5 4 16 16 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 8 7 14 16 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 4 14 16 16 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C16 1 16 4.23171e-15
C15 2 16 7.50427e-16
C14 3 16 7.91113e-16
C13 4 16 3.53148e-14
C12 5 16 1.80046e-15
C11 6 16 1.47638e-14
C10 7 16 1.75794e-14
C8 9 16 1.47638e-14
C7 10 16 1.54677e-14
C6 11 16 1.51158e-14
C3 14 16 1.91094e-14
C2 15 16 1.51158e-14
C1 16 16 3.35293e-15
.ends noa2a2a23_x4

