* Spice description of na3_x4
* Spice driver version -935764197
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:17

* INTERF i0 i1 i2 nq vdd vss 


.subckt na3_x4 8 3 7 5 1 6 
* NET 1 = vdd
* NET 3 = i1
* NET 5 = nq
* NET 6 = vss
* NET 7 = i2
* NET 8 = i0
Xtr_00012 1 2 5 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 5 2 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 1 3 10 1 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Xtr_00009 10 7 1 1 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Xtr_00008 1 8 10 1 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Xtr_00007 2 10 1 1 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00006 6 2 5 6 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00005 5 2 6 6 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00004 4 7 9 6 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00003 6 3 4 6 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00002 2 10 6 6 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00001 9 8 10 6 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
C10 1 6 2.08674e-15
C9 2 6 3.73407e-14
C8 3 6 1.46876e-14
C6 5 6 1.71774e-15
C5 6 6 2.43438e-15
C4 7 6 1.46876e-14
C3 8 6 1.61992e-14
C1 10 6 1.76796e-14
.ends na3_x4

