* Spice description of nmx3_x1
* Spice driver version 658792219
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:20

* INTERF cmd0 cmd1 i0 i1 i2 nq vdd vss 


.subckt nmx3_x1 9 15 6 10 12 14 5 16 
* NET 5 = vdd
* NET 6 = i0
* NET 9 = cmd0
* NET 10 = i1
* NET 12 = i2
* NET 14 = nq
* NET 15 = cmd1
* NET 16 = vss
Xtr_00018 3 12 4 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00017 14 15 3 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00016 5 8 4 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00015 4 10 2 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00014 17 15 5 5 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00013 2 17 14 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00012 1 9 5 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00011 14 6 1 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00010 5 9 8 5 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00009 13 12 18 16 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00008 14 17 13 16 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00007 11 15 14 16 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00006 18 10 11 16 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00005 7 8 16 16 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00004 17 15 16 16 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Xtr_00003 16 9 8 16 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Xtr_00002 14 6 7 16 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00001 16 9 18 16 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
C15 4 16 8.03731e-16
C14 5 16 3.45557e-15
C13 6 16 2.20034e-14
C11 8 16 3.07436e-14
C10 9 16 4.6641e-14
C9 10 16 2.88137e-14
C7 12 16 2.36579e-14
C5 14 16 3.48588e-15
C4 15 16 4.83739e-14
C3 16 16 3.28831e-15
C2 17 16 2.23881e-14
C1 18 16 7.48589e-16
.ends nmx3_x1

