* Spice description of oa2a2a2a24_x4
* Spice driver version -1199456485
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:30

* INTERF i0 i1 i2 i3 i4 i5 i6 i7 q vdd vss 


.subckt oa2a2a2a24_x4 6 5 9 10 12 13 16 17 7 1 19 
* NET 1 = vdd
* NET 5 = i1
* NET 6 = i0
* NET 7 = q
* NET 9 = i2
* NET 10 = i3
* NET 12 = i4
* NET 13 = i5
* NET 16 = i6
* NET 17 = i7
* NET 19 = vss
Xtr_00020 2 5 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00019 1 6 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00018 7 14 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00017 1 14 7 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00016 3 9 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00015 2 10 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00014 3 12 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 4 13 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 4 16 14 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 14 17 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 8 5 14 19 sg13_lv_nmos L=0.13U W=1.67U AS=0.4008P AD=0.4008P PS=3.82U PD=3.82U 
Xtr_00009 19 6 8 19 sg13_lv_nmos L=0.13U W=1.67U AS=0.4008P AD=0.4008P PS=3.82U PD=3.82U 
Xtr_00008 7 14 19 19 sg13_lv_nmos L=0.13U W=1.67U AS=0.4008P AD=0.4008P PS=3.82U PD=3.82U 
Xtr_00007 19 14 7 19 sg13_lv_nmos L=0.13U W=1.67U AS=0.4008P AD=0.4008P PS=3.82U PD=3.82U 
Xtr_00006 19 9 11 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 11 10 14 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 14 12 15 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 15 13 19 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 14 16 18 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 18 17 19 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C19 1 19 4.32693e-15
C18 2 19 7.65866e-16
C17 3 19 1.00274e-15
C16 4 19 1.05788e-15
C15 5 19 1.44119e-14
C14 6 19 1.44119e-14
C13 7 19 1.95175e-15
C11 9 19 1.47638e-14
C10 10 19 1.47638e-14
C8 12 19 1.51158e-14
C7 13 19 1.51158e-14
C6 14 19 3.59233e-14
C4 16 19 1.47638e-14
C3 17 19 1.53915e-14
C1 19 19 3.40924e-15
.ends oa2a2a2a24_x4

