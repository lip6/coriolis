* Spice description of a2_x2
* Spice driver version 753875880
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:30

* INTERF i0 i1 q vdd vss 


.subckt a2_x2 1 2 4 3 7 
* NET 1 = i0
* NET 2 = i1
* NET 3 = vdd
* NET 4 = q
* NET 7 = vss
Mtr_00006 4 5 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 5 1 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00004 3 2 5 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 7 5 4 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 6 2 5 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 7 1 6 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C7 1 7 8.37957e-16
C6 2 7 1.09511e-15
C5 3 7 1.46192e-15
C4 4 7 1.22684e-15
C3 5 7 1.81273e-15
C1 7 7 1.42442e-15
.ends a2_x2

