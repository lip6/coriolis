* Spice description of no3_x4
* Spice driver version 57265064
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:00

* INTERF i0 i1 i2 nq vdd vss 


.subckt no3_x4 1 3 2 8 7 9 
* NET 1 = i0
* NET 2 = i2
* NET 3 = i1
* NET 7 = vdd
* NET 8 = nq
* NET 9 = vss
Mtr_00012 7 10 4 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00011 5 1 10 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00010 7 2 6 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00009 6 3 5 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00008 8 4 7 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00007 7 4 8 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00006 4 10 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00005 10 1 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00004 9 4 8 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 8 4 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 10 2 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00001 9 3 10 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
C10 1 9 8.17567e-16
C9 2 9 8.17567e-16
C8 3 9 9.24715e-16
C7 4 9 1.99373e-15
C4 7 9 2.68231e-15
C3 8 9 1.22684e-15
C2 9 9 2.59659e-15
C1 10 9 3.71378e-15
.ends no3_x4

