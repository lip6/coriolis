* Spice description of ts_x4
* Spice driver version -934093029
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:33

* INTERF cmd i q vdd vss 


.subckt ts_x4 4 3 8 1 7 
* NET 1 = vdd
* NET 3 = i
* NET 4 = cmd
* NET 5 = 4
* NET 7 = vss
* NET 8 = q
Xtr_00012 8 2 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 1 2 8 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 5 4 1 1 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00009 1 4 2 1 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00008 2 5 6 1 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00007 2 3 1 1 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00006 6 3 7 7 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00005 8 6 7 7 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 7 6 8 7 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 5 4 7 7 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 7 5 6 7 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 2 4 6 7 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C8 1 7 3.18881e-15
C7 2 7 4.01796e-14
C6 3 7 1.54884e-14
C5 4 7 5.58087e-14
C4 5 7 2.39072e-14
C3 6 7 3.08055e-14
C2 7 7 2.80048e-15
C1 8 7 1.99345e-15
.ends ts_x4

