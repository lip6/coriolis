* Spice description of oa3ao322_x2
* Spice driver version -1912381669
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:31

* INTERF i0 i1 i2 i3 i4 i5 i6 q vdd vss 


.subckt oa3ao322_x2 12 11 10 7 5 6 8 17 4 16 
* NET 4 = vdd
* NET 5 = i4
* NET 6 = i5
* NET 7 = i3
* NET 8 = i6
* NET 10 = i2
* NET 11 = i1
* NET 12 = i0
* NET 15 = 4
* NET 16 = vss
* NET 17 = q
Xtr_00016 2 7 15 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00015 1 5 2 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00014 3 6 1 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00013 15 8 3 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00012 3 12 4 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00011 4 11 3 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00010 3 10 4 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00009 4 15 17 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 16 7 9 16 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Xtr_00007 9 5 16 16 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Xtr_00006 16 6 9 16 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Xtr_00005 9 8 15 16 sg13_lv_nmos L=0.13U W=1.59U AS=0.3816P AD=0.3816P PS=3.67U PD=3.67U 
Xtr_00004 15 10 13 16 sg13_lv_nmos L=0.13U W=1.22U AS=0.2928P AD=0.2928P PS=2.92U PD=2.92U 
Xtr_00003 13 11 14 16 sg13_lv_nmos L=0.13U W=1.22U AS=0.2928P AD=0.2928P PS=2.92U PD=2.92U 
Xtr_00002 16 15 17 16 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Xtr_00001 14 12 16 16 sg13_lv_nmos L=0.13U W=1.22U AS=0.2928P AD=0.2928P PS=2.92U PD=2.92U 
C15 3 16 1.16332e-15
C14 4 16 2.96417e-15
C13 5 16 1.53915e-14
C12 6 16 1.53915e-14
C11 7 16 1.53915e-14
C10 8 16 1.68755e-14
C9 9 16 6.11902e-16
C8 10 16 1.40599e-14
C7 11 16 1.46876e-14
C6 12 16 1.53915e-14
C3 15 16 1.92872e-14
C2 16 16 2.891e-15
C1 17 16 1.99345e-15
.ends oa3ao322_x2

