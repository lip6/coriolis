* Spice description of nmx2_x4
* Spice driver version -119070949
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:20

* INTERF cmd i0 i1 nq vdd vss 


.subckt nmx2_x4 10 11 6 4 3 13 
* NET 3 = vdd
* NET 4 = nq
* NET 6 = i1
* NET 10 = cmd
* NET 11 = i0
* NET 13 = vss
Xtr_00016 3 5 4 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00015 4 5 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00014 5 8 3 3 sg13_lv_pmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Xtr_00013 3 6 2 3 sg13_lv_pmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Xtr_00012 2 12 8 3 sg13_lv_pmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Xtr_00011 8 10 1 3 sg13_lv_pmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Xtr_00010 1 11 3 3 sg13_lv_pmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Xtr_00009 3 10 12 3 sg13_lv_pmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Xtr_00008 13 5 4 13 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00007 4 5 13 13 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00006 5 8 13 13 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Xtr_00005 13 6 9 13 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Xtr_00004 9 10 8 13 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Xtr_00003 8 12 7 13 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Xtr_00002 13 10 12 13 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Xtr_00001 7 11 13 13 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
C11 3 13 4.03259e-15
C10 4 13 1.99345e-15
C9 5 13 3.60063e-14
C8 6 13 1.83395e-14
C6 8 13 3.066e-14
C4 10 13 5.26214e-14
C3 11 13 1.82277e-14
C2 12 13 1.58286e-14
C1 13 13 3.25593e-15
.ends nmx2_x4

