* Spice description of one_x0
* Spice driver version 1861938971
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:32

* INTERF q vdd vss 


.subckt one_x0 2 1 3 
* NET 1 = vdd
* NET 2 = q
* NET 3 = vss
Xtr_00001 2 3 1 1 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
C3 1 3 1.33045e-15
C2 2 3 1.88083e-15
C1 3 3 1.14082e-14
.ends one_x0

