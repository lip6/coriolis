* Spice description of nxr2_x1
* Spice driver version 838659867
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:26

* INTERF i0 i1 nq vdd vss 


.subckt nxr2_x1 8 3 7 2 9 
* NET 2 = vdd
* NET 3 = i1
* NET 7 = nq
* NET 8 = i0
* NET 9 = vss
Xtr_00012 4 3 2 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00011 2 4 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 1 10 7 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 7 3 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 1 8 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 2 8 10 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00006 4 3 9 9 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00005 9 3 6 9 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 6 10 7 9 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 7 4 5 9 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 9 8 10 9 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 5 8 9 9 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C10 1 9 8.63047e-16
C9 2 9 2.08674e-15
C8 3 9 3.12373e-14
C7 4 9 2.7614e-14
C4 7 9 1.91539e-15
C3 8 9 2.69501e-14
C2 9 9 2.08674e-15
C1 10 9 2.86016e-14
.ends nxr2_x1

