* Spice description of noa22_x4
* Spice driver version -1923674341
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:22

* INTERF i0 i1 i2 nq vdd vss 


.subckt noa22_x4 4 7 8 3 2 10 
* NET 2 = vdd
* NET 3 = nq
* NET 4 = i0
* NET 7 = i1
* NET 8 = i2
* NET 10 = vss
Xtr_00012 2 6 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 2 9 6 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00010 1 4 9 2 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00009 9 7 1 2 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00008 1 8 2 2 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00007 3 6 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 10 6 3 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 10 9 6 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00004 10 4 5 10 sg13_lv_nmos L=0.13U W=1.14U AS=0.2736P AD=0.2736P PS=2.77U PD=2.77U 
Xtr_00003 5 7 9 10 sg13_lv_nmos L=0.13U W=1.14U AS=0.2736P AD=0.2736P PS=2.77U PD=2.77U 
Xtr_00002 9 8 10 10 sg13_lv_nmos L=0.13U W=1.14U AS=0.2736P AD=0.2736P PS=2.77U PD=2.77U 
Xtr_00001 3 6 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C10 1 10 4.31523e-16
C9 2 10 3.40524e-15
C8 3 10 2.02102e-15
C7 4 10 2.76544e-14
C5 6 10 4.3149e-14
C4 7 10 2.70057e-14
C3 8 10 1.8559e-14
C2 9 10 2.07676e-14
C1 10 10 2.93362e-15
.ends noa22_x4

