* Spice description of tie_x0
* Spice driver version 911571880
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:34

* INTERF vdd vss 


.subckt tie_x0 1 2 
* NET 1 = vdd
* NET 2 = vss
C2 1 2 2.89745e-16
C1 2 2 2.89745e-16
.ends tie_x0

