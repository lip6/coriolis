* Spice description of o4_x2
* Spice driver version 139452187
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:28

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt o4_x2 7 8 6 9 5 2 11 
* NET 2 = vdd
* NET 5 = q
* NET 6 = i2
* NET 7 = i0
* NET 8 = i1
* NET 9 = i3
* NET 11 = vss
Xtr_00010 2 6 3 2 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00009 3 7 1 2 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00008 1 8 4 2 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00007 4 9 10 2 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00006 5 10 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00005 11 6 10 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00004 10 7 11 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00003 11 8 10 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 10 9 11 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 5 10 11 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C10 2 11 1.79971e-15
C7 5 11 1.99345e-15
C6 6 11 1.51158e-14
C5 7 11 1.58197e-14
C4 8 11 1.98407e-14
C3 9 11 2.01926e-14
C2 10 11 2.10053e-14
C1 11 11 2.28515e-15
.ends o4_x2

