* Spice description of noa22_x4
* Spice driver version -935949400
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:03

* INTERF i0 i1 i2 nq vdd vss 


.subckt noa22_x4 3 5 4 8 6 10 
* NET 3 = i0
* NET 4 = i2
* NET 5 = i1
* NET 6 = vdd
* NET 8 = nq
* NET 10 = vss
Mtr_00012 6 7 2 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00011 6 4 1 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00010 7 3 1 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00009 1 5 7 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00008 6 2 8 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00007 8 2 6 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00006 2 7 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00005 7 4 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00004 9 5 7 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00003 10 3 9 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00002 10 2 8 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 8 2 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C10 1 10 4.33949e-16
C9 2 10 1.99373e-15
C8 3 10 1.16072e-15
C7 4 10 9.46424e-16
C6 5 10 1.19053e-15
C5 6 10 2.68231e-15
C4 7 10 2.53515e-15
C3 8 10 1.22684e-15
C1 10 10 2.59659e-15
.ends noa22_x4

