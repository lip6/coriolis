* Spice description of inv_x4
* Spice driver version 1333574568
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:43

* INTERF i nq vdd vss 


.subckt inv_x4 1 4 2 3 
* NET 1 = i
* NET 2 = vdd
* NET 3 = vss
* NET 4 = nq
Mtr_00004 2 1 4 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00003 4 1 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00002 4 1 3 3 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 3 1 4 3 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C4 1 3 1.13955e-15
C3 2 3 1.99927e-15
C2 3 3 1.50103e-15
C1 4 3 1.22684e-15
.ends inv_x4

