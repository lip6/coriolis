* Spice description of a4_x2
* Spice driver version 354148123
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:11

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt a4_x2 8 9 4 3 2 1 11 
* NET 1 = vdd
* NET 2 = q
* NET 3 = i3
* NET 4 = i2
* NET 8 = i0
* NET 9 = i1
* NET 11 = vss
Xtr_00010 2 7 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 1 3 7 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00008 7 4 1 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00007 7 8 1 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00006 1 9 7 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00005 7 3 6 11 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00004 2 7 11 11 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Xtr_00003 6 4 5 11 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00002 10 8 11 11 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00001 5 9 10 11 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
C11 1 11 2.61062e-15
C10 2 11 1.93831e-15
C9 3 11 2.01651e-14
C8 4 11 1.57159e-14
C5 7 11 1.80612e-14
C4 8 11 1.47363e-14
C3 9 11 1.5012e-14
C1 11 11 2.06464e-15
.ends a4_x2

