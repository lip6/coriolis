* Spice description of oa2a22_x4
* Spice driver version -1049809125
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:29

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt oa2a22_x4 9 8 4 5 3 2 11 
* NET 2 = vdd
* NET 3 = q
* NET 4 = i2
* NET 5 = i3
* NET 8 = i1
* NET 9 = i0
* NET 11 = vss
Xtr_00012 2 4 1 2 sg13_lv_pmos L=0.13U W=1.59U AS=0.3816P AD=0.3816P PS=3.67U PD=3.67U 
Xtr_00011 1 5 2 2 sg13_lv_pmos L=0.13U W=1.59U AS=0.3816P AD=0.3816P PS=3.67U PD=3.67U 
Xtr_00010 1 8 7 2 sg13_lv_pmos L=0.13U W=1.59U AS=0.3816P AD=0.3816P PS=3.67U PD=3.67U 
Xtr_00009 7 9 1 2 sg13_lv_pmos L=0.13U W=1.59U AS=0.3816P AD=0.3816P PS=3.67U PD=3.67U 
Xtr_00008 3 7 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 2 7 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 6 4 7 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00005 7 8 10 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00004 10 9 11 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00003 3 7 11 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 11 7 3 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 11 5 6 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C11 1 11 8.73826e-16
C10 2 11 3.58371e-15
C9 3 11 1.99345e-15
C8 4 11 2.45421e-14
C7 5 11 2.52459e-14
C5 7 11 4.07614e-14
C4 8 11 2.13745e-14
C3 9 11 2.10226e-14
C1 11 11 3.10676e-15
.ends oa2a22_x4

