* Spice description of ao22_x4
* Spice driver version -49991909
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:12

* INTERF i0 i1 i2 q vdd vss 


.subckt ao22_x4 7 4 5 3 2 6 
* NET 2 = vdd
* NET 3 = q
* NET 4 = i1
* NET 5 = i2
* NET 6 = vss
* NET 7 = i0
Xtr_00010 2 8 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 3 8 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 2 5 8 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00007 8 4 1 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00006 1 7 2 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00005 9 4 8 6 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00004 8 7 9 6 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00003 6 8 3 6 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00002 3 8 6 6 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00001 6 5 9 6 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
C8 2 6 3.50537e-15
C7 3 6 1.93831e-15
C6 4 6 1.80968e-14
C5 5 6 2.09881e-14
C4 6 6 2.61776e-15
C3 7 6 1.74691e-14
C2 8 6 3.96706e-14
C1 9 6 4.45309e-16
.ends ao22_x4

