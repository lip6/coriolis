* Spice description of noa22_x1
* Spice driver version 1328053160
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:02

* INTERF i0 i1 i2 nq vdd vss 


.subckt noa22_x1 1 3 2 7 4 6 
* NET 1 = i0
* NET 2 = i2
* NET 3 = i1
* NET 4 = vdd
* NET 6 = vss
* NET 7 = nq
Mtr_00006 4 2 5 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 7 1 5 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00004 5 3 7 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00003 6 1 8 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 8 3 7 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 7 2 6 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C8 1 6 8.60287e-16
C7 2 6 9.67435e-16
C6 3 6 9.67435e-16
C5 4 6 1.21548e-15
C4 5 6 6.5896e-16
C3 6 6 1.46192e-15
C2 7 6 1.07148e-15
.ends noa22_x1

