* Spice description of oa3ao322_x4
* Spice driver version -79270117
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:31

* INTERF i0 i1 i2 i3 i4 i5 i6 q vdd vss 


.subckt oa3ao322_x4 12 11 9 8 5 6 7 16 4 17 
* NET 4 = vdd
* NET 5 = i4
* NET 6 = i5
* NET 7 = i6
* NET 8 = i3
* NET 9 = i2
* NET 11 = i1
* NET 12 = i0
* NET 16 = q
* NET 17 = vss
Xtr_00018 1 8 15 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00017 2 5 1 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00016 3 6 2 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00015 15 7 3 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00014 3 9 4 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00013 4 11 3 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00012 3 12 4 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00011 4 15 16 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 16 15 4 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 17 8 10 17 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00008 10 7 15 17 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00007 17 6 10 17 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00006 10 5 17 17 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00005 15 9 13 17 sg13_lv_nmos L=0.13U W=1.22U AS=0.2928P AD=0.2928P PS=2.92U PD=2.92U 
Xtr_00004 13 11 14 17 sg13_lv_nmos L=0.13U W=1.22U AS=0.2928P AD=0.2928P PS=2.92U PD=2.92U 
Xtr_00003 14 12 17 17 sg13_lv_nmos L=0.13U W=1.22U AS=0.2928P AD=0.2928P PS=2.92U PD=2.92U 
Xtr_00002 16 15 17 17 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00001 17 15 16 17 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
C15 3 17 1.20468e-15
C14 4 17 4.17826e-15
C13 5 17 1.67993e-14
C12 6 17 1.71512e-14
C11 7 17 1.47776e-14
C10 8 17 1.8207e-14
C9 9 17 1.8649e-14
C8 10 17 5.28022e-16
C7 11 17 2.45808e-14
C6 12 17 2.49328e-14
C3 15 17 4.18428e-14
C2 16 17 1.99345e-15
C1 17 17 3.62334e-15
.ends oa3ao322_x4

