* Spice description of mx2_x2
* Spice driver version -792630360
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:45

* INTERF cmd i0 i1 q vdd vss 


.subckt mx2_x2 7 5 6 4 3 12 
* NET 3 = vdd
* NET 4 = q
* NET 5 = i0
* NET 6 = i1
* NET 7 = cmd
* NET 12 = vss
Mtr_00012 4 10 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00011 1 6 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00010 9 7 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.02U AS=0.2958P AD=0.2958P PS=2.62U PD=2.62U 
Mtr_00009 3 5 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00008 10 9 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00007 2 7 10 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00006 12 6 11 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00005 4 10 12 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00004 12 7 9 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.54U AS=0.1566P AD=0.1566P PS=1.66U PD=1.66U 
Mtr_00003 11 7 10 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00002 8 5 12 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00001 10 9 8 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
C10 3 12 2.51249e-15
C9 4 12 1.22684e-15
C8 5 12 1.05272e-15
C7 6 12 1.11439e-15
C6 7 12 1.49322e-15
C4 9 12 3.46344e-15
C3 10 12 1.92357e-15
C1 12 12 2.18033e-15
.ends mx2_x2

