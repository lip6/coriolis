* Spice description of oa2a2a2a24_x2
* Spice driver version -293425381
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:30

* INTERF i0 i1 i2 i3 i4 i5 i6 i7 q vdd vss 


.subckt oa2a2a2a24_x2 7 6 9 10 13 14 12 17 5 2 19 
* NET 2 = vdd
* NET 5 = q
* NET 6 = i1
* NET 7 = i0
* NET 9 = i2
* NET 10 = i3
* NET 12 = i6
* NET 13 = i4
* NET 14 = i5
* NET 17 = i7
* NET 19 = vss
Xtr_00018 1 6 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00017 2 7 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00016 16 17 4 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00015 5 16 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00014 4 12 16 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 3 9 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 1 10 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 3 13 4 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 4 14 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 8 6 16 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00008 19 7 8 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00007 18 17 19 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00006 5 16 19 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 16 12 18 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 19 9 11 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 11 10 16 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 16 13 15 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 15 14 19 19 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C19 1 19 8.40703e-16
C18 2 19 3.69579e-15
C17 3 19 1.0009e-15
C16 4 19 1.26767e-15
C15 5 19 1.73337e-15
C14 6 19 1.47638e-14
C13 7 19 1.53915e-14
C11 9 19 1.51158e-14
C10 10 19 1.47638e-14
C8 12 19 2.22545e-14
C7 13 19 1.51158e-14
C6 14 19 1.54677e-14
C4 16 19 2.02548e-14
C3 17 19 1.53915e-14
C1 19 19 3.35293e-15
.ends oa2a2a2a24_x2

