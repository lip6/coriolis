* Spice description of o2_x4
* Spice driver version 1602862875
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:27

* INTERF i0 i1 q vdd vss 


.subckt o2_x4 3 5 4 1 6 
* NET 1 = vdd
* NET 3 = i0
* NET 4 = q
* NET 5 = i1
* NET 6 = vss
Xtr_00009 1 7 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 4 7 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 2 5 7 1 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00006 1 3 2 1 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00005 6 7 4 6 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 4 7 6 6 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 6 3 7 6 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 7 5 6 6 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 6 3 7 6 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C7 1 6 2.26478e-15
C5 3 6 1.72387e-14
C4 4 6 1.99345e-15
C3 5 6 1.96148e-14
C2 6 6 2.14138e-15
C1 7 6 3.57653e-14
.ends o2_x4

