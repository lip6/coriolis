* Spice description of buf_x2
* Spice driver version 1659420443
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:13

* INTERF i q vdd vss 


.subckt buf_x2 3 2 1 4 
* NET 1 = vdd
* NET 2 = q
* NET 3 = i
* NET 4 = vss
Xtr_00004 2 5 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00003 1 3 5 1 sg13_lv_pmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00002 4 3 5 4 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Xtr_00001 2 5 4 4 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C5 1 4 1.10757e-15
C4 2 4 1.93831e-15
C3 3 4 1.88002e-14
C2 4 4 1.10757e-15
C1 5 4 3.0571e-14
.ends buf_x2

