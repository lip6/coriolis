* Spice description of ao22_x2
* Spice driver version -1352500312
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:36

* INTERF i0 i1 i2 q vdd vss 


.subckt ao22_x2 3 2 4 6 5 8 
* NET 2 = i1
* NET 3 = i0
* NET 4 = i2
* NET 5 = vdd
* NET 6 = q
* NET 8 = vss
Mtr_00008 1 2 7 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00007 5 3 1 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00006 7 4 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00005 5 7 6 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00004 8 4 9 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00003 9 2 7 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00002 7 3 9 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00001 6 7 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C8 2 8 1.03326e-15
C7 3 8 1.15106e-15
C6 4 8 1.32091e-15
C5 5 8 1.63174e-15
C4 6 8 1.22684e-15
C3 7 8 1.82821e-15
C2 8 8 1.3853e-15
C1 9 8 4.33949e-16
.ends ao22_x2

