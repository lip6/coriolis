* Spice description of nao2o22_x4
* Spice driver version 2054246171
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:19

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt nao2o22_x4 10 7 6 8 4 3 9 
* NET 3 = vdd
* NET 4 = nq
* NET 6 = i2
* NET 7 = i1
* NET 8 = i3
* NET 9 = vss
* NET 10 = i0
Xtr_00014 1 8 11 3 sg13_lv_pmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
Xtr_00013 3 6 1 3 sg13_lv_pmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
Xtr_00012 11 7 2 3 sg13_lv_pmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
Xtr_00011 4 5 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 3 5 4 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 2 10 3 3 sg13_lv_pmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
Xtr_00008 3 11 5 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00007 12 6 9 9 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00006 4 5 9 9 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 9 5 4 9 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 12 7 11 9 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00003 11 10 12 9 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00002 9 11 5 9 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 9 8 12 9 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
C10 3 9 3.67183e-15
C9 4 9 1.99345e-15
C8 5 9 3.99639e-14
C7 6 9 2.71959e-14
C6 7 9 2.43397e-14
C5 8 9 2.35092e-14
C4 9 9 3.25477e-15
C3 10 9 1.8559e-14
C2 11 9 2.18104e-14
C1 12 9 8.18684e-16
.ends nao2o22_x4

