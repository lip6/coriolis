* Spice description of noa2a22_x1
* Spice driver version -496750821
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:22

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt noa2a22_x1 8 7 4 3 6 1 10 
* NET 1 = vdd
* NET 3 = i3
* NET 4 = i2
* NET 6 = nq
* NET 7 = i1
* NET 8 = i0
* NET 10 = vss
Xtr_00008 2 7 6 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 6 8 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 1 3 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00005 2 4 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00004 6 7 9 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 9 8 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 5 3 6 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 10 4 5 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C10 1 10 1.569e-15
C9 2 10 8.6004e-16
C8 3 10 1.53152e-14
C7 4 10 1.6723e-14
C5 6 10 1.89763e-15
C4 7 10 1.50395e-14
C3 8 10 1.50395e-14
C1 10 10 1.62531e-15
.ends noa2a22_x1

