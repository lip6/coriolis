* Spice description of oa2ao222_x2
* Spice driver version 154930971
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:30

* INTERF i0 i1 i2 i3 i4 q vdd vss 


.subckt oa2ao222_x2 11 10 6 4 7 5 3 13 
* NET 3 = vdd
* NET 4 = i3
* NET 5 = q
* NET 6 = i2
* NET 7 = i4
* NET 10 = i1
* NET 11 = i0
* NET 13 = vss
Xtr_00012 2 4 1 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 1 6 8 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 2 10 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 3 11 2 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 8 7 2 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 5 8 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 9 4 13 13 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Xtr_00005 13 6 9 13 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Xtr_00004 12 11 13 13 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Xtr_00003 8 10 12 13 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Xtr_00002 9 7 8 13 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Xtr_00001 5 8 13 13 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
C12 2 13 9.28968e-16
C11 3 13 2.49967e-15
C10 4 13 1.4838e-14
C9 5 13 2.04976e-15
C8 6 13 1.79701e-14
C7 7 13 1.50299e-14
C6 8 13 1.20682e-14
C5 9 13 4.45309e-16
C4 10 13 1.60095e-14
C3 11 13 1.59333e-14
C1 13 13 2.69383e-15
.ends oa2ao222_x2

