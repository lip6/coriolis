* Spice description of a4_x4
* Spice driver version 1435143080
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:34

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt a4_x4 4 5 1 2 11 7 8 
* NET 1 = i2
* NET 2 = i3
* NET 4 = i0
* NET 5 = i1
* NET 7 = vdd
* NET 8 = vss
* NET 11 = q
Mtr_00012 11 6 7 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00011 7 6 11 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00010 7 5 6 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00009 7 2 6 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00008 6 1 7 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00007 6 4 7 7 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00006 8 6 11 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00005 11 6 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00004 8 4 10 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 3 2 6 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 9 1 3 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 10 5 9 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C11 1 8 1.04216e-15
C10 2 8 1.09479e-15
C8 4 8 1.04216e-15
C7 5 8 9.82537e-16
C6 6 8 2.76982e-15
C5 7 8 3.71629e-15
C4 8 8 2.55909e-15
C1 11 8 1.22684e-15
.ends a4_x4

