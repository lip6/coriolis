* Spice description of noa2a2a2a24_x1
* Spice driver version -970170597
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:24

* INTERF i0 i1 i2 i3 i4 i5 i6 i7 nq vdd vss 


.subckt noa2a2a2a24_x1 6 5 8 9 11 12 13 16 15 1 18 
* NET 1 = vdd
* NET 5 = i1
* NET 6 = i0
* NET 8 = i2
* NET 9 = i3
* NET 11 = i4
* NET 12 = i5
* NET 13 = i6
* NET 15 = nq
* NET 16 = i7
* NET 18 = vss
Xtr_00016 2 5 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00015 1 6 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00014 2 9 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 3 8 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 3 11 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 4 12 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 4 13 15 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 15 16 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 7 5 15 18 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00007 18 6 7 18 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00006 18 8 10 18 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00005 10 9 15 18 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00004 15 11 14 18 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00003 14 12 18 18 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00002 15 13 17 18 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00001 17 16 18 18 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
C18 1 18 2.93601e-15
C17 2 18 7.8987e-16
C16 3 18 1.0009e-15
C15 4 18 1.26767e-15
C14 5 18 1.51158e-14
C13 6 18 1.50395e-14
C11 8 18 2.20688e-14
C10 9 18 2.17169e-14
C8 11 18 2.17169e-14
C7 12 18 2.17169e-14
C6 13 18 2.04337e-14
C4 15 18 2.67991e-15
C3 16 18 2.20064e-14
C1 18 18 3.03119e-15
.ends noa2a2a2a24_x1

