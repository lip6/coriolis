* Spice description of nao22_x4
* Spice driver version 1184426920
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:53

* INTERF i0 i1 i2 nq vdd vss 


.subckt nao22_x4 3 5 4 7 6 9 
* NET 3 = i0
* NET 4 = i2
* NET 5 = i1
* NET 6 = vdd
* NET 7 = nq
* NET 9 = vss
Mtr_00012 6 8 2 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00011 6 4 8 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00010 1 3 6 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00009 8 5 1 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00008 6 2 7 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00007 7 2 6 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00006 2 8 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00005 10 4 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00004 8 5 10 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00003 10 3 8 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00002 9 2 7 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 7 2 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C9 2 9 1.99373e-15
C8 3 9 1.16072e-15
C7 4 9 9.46424e-16
C6 5 9 1.19053e-15
C5 6 9 2.92875e-15
C4 7 9 1.22684e-15
C3 8 9 2.53515e-15
C2 9 9 2.35015e-15
C1 10 9 8.08967e-16
.ends nao22_x4

