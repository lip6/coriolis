* Spice description of no4_x1
* Spice driver version 145178395
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:21

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt no4_x1 7 8 6 5 9 1 10 
* NET 1 = vdd
* NET 5 = i3
* NET 6 = i2
* NET 7 = i0
* NET 8 = i1
* NET 9 = nq
* NET 10 = vss
Xtr_00008 3 6 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 2 7 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 4 8 9 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00005 1 5 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00004 10 5 9 10 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Xtr_00003 9 6 10 10 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Xtr_00002 10 7 9 10 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Xtr_00001 9 8 10 10 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
C10 1 10 1.569e-15
C6 5 10 2.13371e-14
C5 6 10 1.9251e-14
C4 7 10 2.11354e-14
C3 8 10 1.98531e-14
C2 9 10 2.56699e-15
C1 10 10 2.08691e-15
.ends no4_x1

