* Spice description of noa2a2a23_x4
* Spice driver version 261217192
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:06

* INTERF i0 i1 i2 i3 i4 i5 nq vdd vss 


.subckt noa2a2a23_x4 9 12 10 11 4 5 3 6 16 
* NET 3 = nq
* NET 4 = i4
* NET 5 = i5
* NET 6 = vdd
* NET 9 = i0
* NET 10 = i2
* NET 11 = i3
* NET 12 = i1
* NET 16 = vss
Mtr_00018 2 11 1 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00017 1 10 2 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00016 1 12 14 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00015 6 4 2 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00014 2 5 6 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00013 14 9 1 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00012 7 14 6 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00011 3 7 6 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00010 6 7 3 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00009 8 4 16 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00008 13 10 16 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00007 14 11 13 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00006 15 12 14 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00005 16 9 15 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00004 14 5 8 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
Mtr_00003 16 7 3 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 3 7 16 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 16 14 7 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
C16 1 16 1.20006e-15
C15 2 16 7.87538e-16
C14 3 16 1.22684e-15
C13 4 16 9.46424e-16
C12 5 16 9.19745e-16
C11 6 16 4.90131e-15
C10 7 16 1.8253e-15
C8 9 16 1.07871e-15
C7 10 16 9.46424e-16
C6 11 16 8.39275e-16
C5 12 16 1.05357e-15
C3 14 16 3.19052e-15
C1 16 16 4.31735e-15
.ends noa2a2a23_x4

