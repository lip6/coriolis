* Spice description of oa22_x2
* Spice driver version 1876659995
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:28

* INTERF i0 i1 i2 q vdd vss 


.subckt oa22_x2 6 7 3 4 2 9 
* NET 2 = vdd
* NET 3 = i2
* NET 4 = q
* NET 6 = i0
* NET 7 = i1
* NET 9 = vss
Xtr_00008 4 5 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 1 7 5 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00006 2 3 1 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00005 5 6 1 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00004 4 5 9 9 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 9 3 5 9 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 5 7 8 9 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 8 6 9 9 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C9 1 9 6.68882e-16
C8 2 9 1.569e-15
C7 3 9 1.71681e-14
C6 4 9 1.99345e-15
C5 5 9 2.0875e-14
C4 6 9 2.27823e-14
C3 7 9 1.54884e-14
C1 9 9 1.62531e-15
.ends oa22_x2

