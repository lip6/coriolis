* Spice description of noa2a22_x1
* Spice driver version 687975336
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:03

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt noa2a22_x1 4 3 2 1 8 6 9 
* NET 1 = i3
* NET 2 = i2
* NET 3 = i1
* NET 4 = i0
* NET 6 = vdd
* NET 8 = nq
* NET 9 = vss
Mtr_00008 6 1 5 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00007 5 2 6 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00006 5 3 8 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 8 4 5 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00004 7 2 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 8 1 7 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 10 3 8 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 9 4 10 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C10 1 9 9.67435e-16
C9 2 9 8.038e-16
C8 3 9 8.60287e-16
C7 4 9 8.85424e-16
C6 5 9 1.484e-15
C5 6 9 1.3853e-15
C3 8 9 1.24827e-15
C2 9 9 1.63174e-15
.ends noa2a22_x1

