* Spice description of mx2_x2
* Spice driver version -1308258533
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:15

* INTERF cmd i0 i1 q vdd vss 


.subckt mx2_x2 9 10 4 5 3 11 
* NET 3 = vdd
* NET 4 = i1
* NET 5 = q
* NET 9 = cmd
* NET 10 = i0
* NET 11 = vss
Xtr_00012 7 9 2 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00011 1 12 7 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00010 3 4 1 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00009 3 9 12 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00008 2 10 3 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00007 5 7 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 11 4 8 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00005 8 9 7 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00004 7 12 6 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00003 6 10 11 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 11 9 12 11 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 5 7 11 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C10 3 11 2.28632e-15
C9 4 11 1.80023e-14
C8 5 11 1.93831e-15
C6 7 11 2.45636e-14
C4 9 11 6.01647e-14
C3 10 11 2.00085e-14
C2 11 11 2.08674e-15
C1 12 11 1.82808e-14
.ends mx2_x2

