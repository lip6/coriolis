* Spice description of noa3ao322_x4
* Spice driver version 939536155
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:25

* INTERF i0 i1 i2 i3 i4 i5 i6 nq vdd vss 


.subckt noa3ao322_x4 13 10 8 6 7 5 9 15 4 18 
* NET 4 = vdd
* NET 5 = i5
* NET 6 = i3
* NET 7 = i4
* NET 8 = i2
* NET 9 = i6
* NET 10 = i1
* NET 13 = i0
* NET 15 = nq
* NET 18 = vss
Xtr_00020 3 13 4 4 sg13_lv_pmos L=0.13U W=1.67U AS=0.4008P AD=0.4008P PS=3.82U PD=3.82U 
Xtr_00019 16 9 3 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00018 3 8 4 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00017 1 6 16 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00016 2 7 1 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00015 3 5 2 4 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00014 4 10 3 4 sg13_lv_pmos L=0.13U W=1.67U AS=0.4008P AD=0.4008P PS=3.82U PD=3.82U 
Xtr_00013 15 17 4 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 4 17 15 4 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 4 16 17 4 sg13_lv_pmos L=0.13U W=1.82U AS=0.4368P AD=0.4368P PS=4.12U PD=4.12U 
Xtr_00010 16 8 12 18 sg13_lv_nmos L=0.13U W=1.22U AS=0.2928P AD=0.2928P PS=2.92U PD=2.92U 
Xtr_00009 14 13 18 18 sg13_lv_nmos L=0.13U W=1.22U AS=0.2928P AD=0.2928P PS=2.92U PD=2.92U 
Xtr_00008 11 9 16 18 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00007 18 6 11 18 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00006 11 7 18 18 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00005 18 5 11 18 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00004 12 10 14 18 sg13_lv_nmos L=0.13U W=1.22U AS=0.2928P AD=0.2928P PS=2.92U PD=2.92U 
Xtr_00003 15 17 18 18 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00002 18 17 15 18 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00001 18 16 17 18 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
C16 3 18 1.14954e-15
C15 4 18 4.15369e-15
C14 5 18 1.39837e-14
C13 6 18 1.46876e-14
C12 7 18 1.43356e-14
C11 8 18 1.3708e-14
C10 9 18 1.51158e-14
C9 10 18 1.57434e-14
C8 11 18 5.28022e-16
C6 13 18 1.57434e-14
C4 15 18 1.93714e-15
C3 16 18 2.50312e-14
C2 17 18 2.64316e-14
C1 18 18 3.85405e-15
.ends noa3ao322_x4

