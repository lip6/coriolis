* Spice description of a4_x2
* Spice driver version 22121384
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:34

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt a4_x2 5 2 3 1 7 6 8 
* NET 1 = i3
* NET 2 = i1
* NET 3 = i2
* NET 5 = i0
* NET 6 = vdd
* NET 7 = q
* NET 8 = vss
Mtr_00010 4 5 6 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00009 7 4 6 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00008 6 1 4 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00007 4 3 6 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00006 6 2 4 6 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00005 8 5 9 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00004 9 2 10 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 11 1 4 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 10 3 11 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 8 4 7 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C11 1 8 1.09479e-15
C10 2 8 9.82537e-16
C9 3 8 1.04216e-15
C8 4 8 2.57005e-15
C7 5 8 1.04216e-15
C6 6 8 2.75893e-15
C5 7 8 1.22684e-15
C4 8 8 1.93389e-15
.ends a4_x2

