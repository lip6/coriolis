* Spice description of mx3_x2
* Spice driver version -1653113061
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:16

* INTERF cmd0 cmd1 i0 i1 i2 q vdd vss 


.subckt mx3_x2 9 17 7 11 13 6 5 19 
* NET 5 = vdd
* NET 6 = q
* NET 7 = i0
* NET 9 = cmd0
* NET 11 = i1
* NET 13 = i2
* NET 17 = cmd1
* NET 19 = vss
Xtr_00020 4 13 3 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00019 6 16 5 5 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00018 5 9 10 5 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00017 16 17 4 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00016 2 18 16 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00015 3 11 2 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00014 5 10 3 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00013 1 9 5 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00012 16 7 1 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00011 18 17 5 5 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00010 15 13 14 19 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00009 19 9 10 19 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Xtr_00008 6 16 19 19 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Xtr_00007 16 18 15 19 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00006 12 17 16 19 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00005 14 11 12 19 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00004 8 10 19 19 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00003 18 17 19 19 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Xtr_00002 16 7 8 19 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00001 19 9 14 19 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
C17 3 19 7.34803e-16
C15 5 19 3.74668e-15
C14 6 19 2.04976e-15
C13 7 19 2.1941e-14
C11 9 19 4.54419e-14
C10 10 19 3.07557e-14
C9 11 19 2.36681e-14
C7 13 19 2.37976e-14
C6 14 19 7.21018e-16
C4 16 19 1.96303e-14
C3 17 19 4.58965e-14
C2 18 19 1.72385e-14
C1 19 19 3.47767e-15
.ends mx3_x2

