* Spice description of nao22_x1
* Spice driver version -520266840
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:52

* INTERF i0 i1 i2 nq vdd vss 


.subckt nao22_x1 1 3 2 7 5 8 
* NET 1 = i0
* NET 2 = i2
* NET 3 = i1
* NET 5 = vdd
* NET 7 = nq
* NET 8 = vss
Mtr_00006 5 2 7 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 4 1 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00004 7 3 4 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00003 6 1 7 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 7 3 6 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 6 2 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C8 1 8 9.67435e-16
C7 2 8 9.67435e-16
C6 3 8 9.67435e-16
C4 5 8 1.46192e-15
C3 6 8 4.33949e-16
C2 7 8 1.24827e-15
C1 8 8 1.21548e-15
.ends nao22_x1

