* Spice description of sff2_x4
* Spice driver version 1979735835
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:33

* INTERF ck cmd i0 i1 q vdd vss 


.subckt sff2_x4 15 21 22 16 7 6 24 
* NET 6 = vdd
* NET 7 = q
* NET 8 = sff_s
* NET 12 = sff_m
* NET 14 = ckr
* NET 15 = ck
* NET 16 = i1
* NET 17 = nckr
* NET 21 = cmd
* NET 22 = i0
* NET 24 = vss
Xtr_00034 3 17 12 6 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00033 12 14 2 6 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00032 7 8 6 6 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00031 1 14 8 6 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00030 8 17 10 6 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00029 6 10 3 6 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00028 6 8 7 6 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00027 10 12 6 6 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00026 19 21 5 6 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00025 4 23 19 6 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00024 6 16 4 6 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00023 6 15 17 6 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00022 6 7 1 6 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00021 5 22 6 6 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00020 6 21 23 6 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00019 14 17 6 6 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00018 2 19 6 6 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00017 12 17 11 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00016 8 14 10 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00015 7 8 24 24 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00014 13 14 12 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00013 10 12 24 24 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Xtr_00012 24 10 13 24 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Xtr_00011 24 8 7 24 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00010 24 7 9 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00009 19 23 20 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00008 20 22 24 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00007 24 21 23 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00006 24 15 17 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00005 14 17 24 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00004 11 19 24 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00003 9 17 8 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 18 21 19 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 24 16 18 24 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C19 6 24 7.22839e-15
C18 7 24 2.26378e-14
C17 8 24 3.39914e-14
C15 10 24 1.74015e-14
C13 12 24 2.35107e-14
C11 14 24 6.87917e-14
C10 15 24 1.85796e-14
C9 16 24 1.33142e-14
C8 17 24 9.65074e-14
C6 19 24 1.38621e-14
C4 21 24 4.67908e-14
C3 22 24 1.68199e-14
C2 23 24 2.03955e-14
C1 24 24 6.56202e-15
.ends sff2_x4

