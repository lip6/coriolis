* Spice description of nmx2_x1
* Spice driver version 1104228123
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:19

* INTERF cmd i0 i1 nq vdd vss 


.subckt nmx2_x1 8 9 4 7 3 10 
* NET 3 = vdd
* NET 4 = i1
* NET 7 = nq
* NET 8 = cmd
* NET 9 = i0
* NET 10 = vss
* NET 11 = q
Xtr_00010 3 4 1 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 7 8 2 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 2 9 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 3 8 11 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00006 1 11 7 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00005 10 4 5 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 7 11 6 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 6 9 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 10 8 11 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 5 8 7 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C9 3 10 1.85602e-15
C8 4 10 1.9138e-14
C5 7 10 1.66327e-15
C4 8 10 4.22155e-14
C3 9 10 1.19689e-14
C2 10 10 1.85602e-15
C1 11 10 1.52849e-14
.ends nmx2_x1

