* Spice description of no2_x4
* Spice driver version -176578789
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:20

* INTERF i0 i1 nq vdd vss 


.subckt no2_x4 5 6 4 1 8 
* NET 1 = vdd
* NET 4 = nq
* NET 5 = i0
* NET 6 = i1
* NET 8 = vss
Xtr_00010 1 5 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 2 6 7 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 1 3 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 4 3 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 3 7 1 1 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00005 8 5 7 8 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00004 7 6 8 8 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00003 4 3 8 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 8 3 4 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 3 7 8 8 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C8 1 8 1.85602e-15
C6 3 8 3.21505e-14
C5 4 8 1.48222e-15
C4 5 8 1.53915e-14
C3 6 8 1.53915e-14
C2 7 8 2.21735e-14
C1 8 8 2.19172e-15
.ends no2_x4

