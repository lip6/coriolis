* Spice description of ao2o22_x4
* Spice driver version 1826103067
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:13

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt ao2o22_x4 9 8 6 5 4 3 7 
* NET 3 = vdd
* NET 4 = q
* NET 5 = i3
* NET 6 = i2
* NET 7 = vss
* NET 8 = i1
* NET 9 = i0
Xtr_00012 3 5 1 3 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00011 3 10 4 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 4 10 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 1 6 10 3 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00008 10 8 2 3 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00007 2 9 3 3 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00006 11 5 7 7 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00005 7 6 11 7 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00004 7 10 4 7 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 4 10 7 7 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 11 8 10 7 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00001 10 9 11 7 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
C9 3 7 3.23798e-15
C8 4 7 1.93831e-15
C7 5 7 2.69505e-14
C6 6 7 2.66081e-14
C5 7 7 2.7382e-15
C4 8 7 1.85314e-14
C3 9 7 1.82557e-14
C2 10 7 4.1784e-14
C1 11 7 7.49757e-16
.ends ao2o22_x4

