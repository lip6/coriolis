* Spice description of oa2a2a23_x2
* Spice driver version 478379803
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:29

* INTERF i0 i1 i2 i3 i4 i5 q vdd vss 


.subckt oa2a2a23_x2 6 5 8 9 12 13 4 2 15 
* NET 2 = vdd
* NET 4 = q
* NET 5 = i1
* NET 6 = i0
* NET 8 = i2
* NET 9 = i3
* NET 12 = i4
* NET 13 = i5
* NET 15 = vss
Xtr_00014 1 5 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 2 6 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 4 11 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 3 8 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 1 9 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 3 12 11 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 11 13 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 7 5 11 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00006 15 6 7 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00005 4 11 15 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 15 8 10 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 10 9 11 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 11 12 14 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 14 13 15 15 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C15 1 15 7.38296e-16
C14 2 15 3.13433e-15
C13 3 15 7.63542e-16
C12 4 15 1.99345e-15
C11 5 15 1.47638e-14
C10 6 15 1.47638e-14
C8 8 15 1.47638e-14
C7 9 15 1.51158e-14
C5 11 15 1.70376e-14
C4 12 15 1.47638e-14
C3 13 15 1.47638e-14
C1 15 15 2.60448e-15
.ends oa2a2a23_x2

