* Spice description of oa2ao222_x4
* Spice driver version -542638309
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:31

* INTERF i0 i1 i2 i3 i4 q vdd vss 


.subckt oa2ao222_x4 11 10 5 6 7 4 2 13 
* NET 2 = vdd
* NET 4 = q
* NET 5 = i2
* NET 6 = i3
* NET 7 = i4
* NET 10 = i1
* NET 11 = i0
* NET 13 = vss
Xtr_00014 2 8 4 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00013 4 8 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 3 6 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 8 7 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 3 10 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 2 11 3 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00008 1 5 8 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 13 8 4 13 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00006 4 8 13 13 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00005 13 5 9 13 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00004 9 6 13 13 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00003 9 7 8 13 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00002 8 10 12 13 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00001 12 11 13 13 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
C12 2 13 3.60538e-15
C11 3 13 9.15182e-16
C10 4 13 2.04976e-15
C9 5 13 1.61058e-14
C8 6 13 2.74006e-14
C7 7 13 1.44119e-14
C6 8 13 3.68461e-14
C5 9 13 4.45309e-16
C4 10 13 1.44119e-14
C3 11 13 1.50395e-14
C1 13 13 3.71516e-15
.ends oa2ao222_x4

