* Spice description of a2_x4
* Spice driver version -1293481048
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:31

* INTERF i0 i1 q vdd vss 


.subckt a2_x4 2 1 5 3 6 
* NET 1 = i1
* NET 2 = i0
* NET 3 = vdd
* NET 5 = q
* NET 6 = vss
Mtr_00008 3 7 5 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00007 5 7 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00006 3 1 7 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00005 7 2 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00004 6 7 5 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 4 1 7 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 6 2 4 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 5 7 6 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C7 1 6 1.09511e-15
C6 2 6 8.37957e-16
C5 3 6 2.41928e-15
C3 5 6 1.22684e-15
C2 6 6 2.04962e-15
C1 7 6 2.08981e-15
.ends a2_x4

