* Spice description of no3_x4
* Spice driver version -686907621
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:21

* INTERF i0 i1 i2 nq vdd vss 


.subckt no3_x4 5 7 8 6 1 10 
* NET 1 = vdd
* NET 5 = i0
* NET 6 = nq
* NET 7 = i1
* NET 8 = i2
* NET 10 = vss
Xtr_00012 1 5 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 2 7 3 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 3 8 9 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00009 4 9 1 1 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00008 1 4 6 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 6 4 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 10 8 9 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00005 4 9 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 6 4 10 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 10 5 9 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 9 7 10 10 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 10 4 6 10 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C10 1 10 2.08674e-15
C7 4 10 3.54006e-14
C6 5 10 1.78551e-14
C5 6 10 1.5562e-15
C4 7 10 1.78551e-14
C3 8 10 1.57434e-14
C2 9 10 2.23053e-14
C1 10 10 2.08674e-15
.ends no3_x4

