* Spice description of nts_x1
* Spice driver version -563840088
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:58:11

* INTERF cmd i nq vdd vss 


.subckt nts_x1 1 2 8 3 6 
* NET 1 = cmd
* NET 2 = i
* NET 3 = vdd
* NET 6 = vss
* NET 8 = nq
Mtr_00006 8 2 4 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00005 4 5 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00004 5 1 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 8 2 7 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 7 1 6 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 6 1 5 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.66U AS=0.1914P AD=0.1914P PS=1.9U PD=1.9U 
C8 1 6 1.10285e-15
C7 2 6 1.18173e-15
C6 3 6 1.36013e-15
C4 5 6 1.30376e-15
C3 6 6 1.21548e-15
C1 8 6 1.22684e-15
.ends nts_x1

