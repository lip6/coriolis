* Spice description of mx3_x4
* Spice driver version 812166939
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:16

* INTERF cmd0 cmd1 i0 i1 i2 q vdd vss 


.subckt mx3_x4 8 16 7 10 12 6 5 18 
* NET 5 = vdd
* NET 6 = q
* NET 7 = i0
* NET 8 = cmd0
* NET 10 = i1
* NET 12 = i2
* NET 16 = cmd1
* NET 18 = vss
Xtr_00022 5 8 9 5 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00021 5 15 6 5 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00020 6 15 5 5 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00019 4 10 3 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00018 15 7 1 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00017 3 19 15 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00016 5 9 4 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00015 1 8 5 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00014 2 12 4 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00013 19 16 5 5 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00012 15 16 2 5 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00011 18 8 9 18 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Xtr_00010 18 15 6 18 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00009 6 15 18 18 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00008 11 9 18 18 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00007 19 16 18 18 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Xtr_00006 14 12 17 18 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00005 15 19 14 18 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00004 13 16 15 18 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00003 17 10 13 18 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00002 15 7 11 18 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Xtr_00001 18 8 17 18 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
C16 4 18 7.7616e-16
C15 5 18 4.67336e-15
C14 6 18 2.2446e-15
C13 7 18 2.3532e-14
C12 8 18 4.89787e-14
C11 9 18 3.20805e-14
C10 10 18 3.18977e-14
C8 12 18 3.25523e-14
C5 15 18 3.5902e-14
C4 16 18 5.02108e-14
C3 17 18 7.48589e-16
C2 18 18 4.19931e-15
C1 19 18 1.93794e-14
.ends mx3_x4

