* Spice description of a3_x2
* Spice driver version 302410664
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2024 at 18:57:32

* INTERF i0 i1 i2 q vdd vss 


.subckt a3_x2 2 1 3 5 4 7 
* NET 1 = i1
* NET 2 = i0
* NET 3 = i2
* NET 4 = vdd
* NET 5 = q
* NET 7 = vss
Mtr_00008 9 3 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00007 5 9 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.7134P AD=0.7134P PS=5.5U PD=5.5U 
Mtr_00006 9 2 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00005 4 1 9 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00004 6 3 9 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00003 7 9 5 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00002 8 1 6 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
Mtr_00001 7 2 8 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.26U AS=0.3654P AD=0.3654P PS=3.1U PD=3.1U 
C9 1 7 9.89144e-16
C8 2 7 8.39136e-16
C7 3 7 9.89143e-16
C6 4 7 1.63174e-15
C5 5 7 1.22684e-15
C3 7 7 1.59424e-15
C1 9 7 2.54251e-15
.ends a3_x2

