* Spice description of buf_x4
* Spice driver version -1111933157
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:14

* INTERF i q vdd vss 


.subckt buf_x4 3 2 1 4 
* NET 1 = vdd
* NET 2 = q
* NET 3 = i
* NET 4 = vss
Xtr_00006 1 5 2 1 sg13_lv_pmos L=0.13U W=2.87U AS=0.6888P AD=0.6888P PS=6.22U PD=6.22U 
Xtr_00005 2 5 1 1 sg13_lv_pmos L=0.13U W=2.87U AS=0.6888P AD=0.6888P PS=6.22U PD=6.22U 
Xtr_00004 1 3 5 1 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00003 4 5 2 4 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00002 2 5 4 4 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00001 4 3 5 4 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C5 1 4 2.02028e-15
C4 2 4 1.93831e-15
C3 3 4 2.05599e-14
C2 4 4 1.63195e-15
C1 5 4 4.69917e-14
.ends buf_x4

