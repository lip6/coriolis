* Spice description of a4_x4
* Spice driver version -233447653
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:11

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt a4_x4 8 9 4 3 2 1 11 
* NET 1 = vdd
* NET 2 = q
* NET 3 = i3
* NET 4 = i2
* NET 8 = i0
* NET 9 = i1
* NET 11 = vss
Xtr_00012 1 7 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 1 3 7 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00010 7 4 1 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00009 1 9 7 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00008 7 8 1 1 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00007 2 7 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 7 3 6 11 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00005 11 7 2 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00004 2 7 11 11 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 6 4 5 11 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00002 10 8 11 11 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00001 5 9 10 11 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
C11 1 11 3.56469e-15
C10 2 11 1.93831e-15
C9 3 11 2.06059e-14
C8 4 11 1.67441e-14
C5 7 11 3.59331e-14
C4 8 11 1.47087e-14
C3 9 11 1.56883e-14
C1 11 11 2.56145e-15
.ends a4_x4

