* Spice description of noa22_x1
* Spice driver version 1120378651
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:22

* INTERF i0 i1 i2 nq vdd vss 


.subckt noa22_x1 6 5 3 4 1 8 
* NET 1 = vdd
* NET 3 = i2
* NET 4 = nq
* NET 5 = i1
* NET 6 = i0
* NET 8 = vss
Xtr_00006 1 3 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00005 2 5 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00004 4 6 2 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00003 8 3 4 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 4 5 7 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 7 6 8 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C8 1 8 1.33828e-15
C7 2 8 6.41311e-16
C6 3 8 2.05182e-14
C5 4 8 1.91482e-15
C4 5 8 1.47638e-14
C3 6 8 1.60954e-14
C1 8 8 1.39459e-15
.ends noa22_x1

