* Spice description of o2_x2
* Spice driver version -524144869
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:26

* INTERF i0 i1 q vdd vss 


.subckt o2_x2 3 5 4 1 7 
* NET 1 = vdd
* NET 3 = i0
* NET 4 = q
* NET 5 = i1
* NET 7 = vss
Xtr_00006 2 5 6 1 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00005 4 6 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00004 1 3 2 1 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Xtr_00003 7 3 6 7 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00002 6 5 7 7 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Xtr_00001 4 6 7 7 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C7 1 7 1.33828e-15
C5 3 7 1.60398e-14
C4 4 7 1.99345e-15
C3 5 7 2.10614e-14
C2 6 7 2.09836e-14
C1 7 7 1.52357e-15
.ends o2_x2

