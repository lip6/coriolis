* Spice description of inv_x8
* Spice driver version -937222373
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:15

* INTERF i nq vdd vss 


.subckt inv_x8 2 4 1 3 
* NET 1 = vdd
* NET 2 = i
* NET 3 = vss
* NET 4 = nq
Xtr_00008 4 2 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00007 1 2 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00006 4 2 1 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00005 1 2 4 1 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00004 4 2 3 3 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00003 3 2 4 3 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 4 2 3 3 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 3 2 4 3 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C4 1 3 2.93299e-15
C3 2 3 8.01992e-14
C2 3 3 2.15634e-15
C1 4 3 3.29763e-15
.ends inv_x8

