* Spice description of nts_x1
* Spice driver version -1531891941
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:25

* INTERF cmd i nq vdd vss 


.subckt nts_x1 5 6 4 2 8 
* NET 2 = vdd
* NET 4 = nq
* NET 5 = cmd
* NET 6 = i
* NET 8 = vss
Xtr_00006 4 3 1 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00005 1 6 2 2 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00004 2 5 3 2 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00003 4 5 7 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00002 7 6 8 8 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Xtr_00001 8 5 3 8 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C7 2 8 2.09702e-15
C6 3 8 1.23468e-14
C5 4 8 1.99345e-15
C4 5 8 3.10765e-14
C3 6 8 1.62948e-14
C1 8 8 1.765e-15
.ends nts_x1

