* Spice description of noa2ao222_x4
* Spice driver version -677781733
* Date ( dd/mm/yyyy hh:mm:ss ): 21/12/2024 at 16:03:24

* INTERF i0 i1 i2 i3 i4 nq vdd vss 


.subckt noa2ao222_x4 10 11 7 5 8 4 3 14 
* NET 3 = vdd
* NET 4 = nq
* NET 5 = i3
* NET 7 = i2
* NET 8 = i4
* NET 10 = i0
* NET 11 = i1
* NET 14 = vss
Xtr_00016 1 7 13 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00015 2 5 1 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00014 2 11 3 3 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00013 3 6 4 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00012 4 6 3 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00011 13 8 2 3 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Xtr_00010 3 10 2 3 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Xtr_00009 3 13 6 3 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00008 9 5 14 14 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Xtr_00007 14 7 9 14 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00006 9 8 13 14 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00005 14 6 4 14 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00004 4 6 14 14 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Xtr_00003 12 10 14 14 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00002 13 11 12 14 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Xtr_00001 14 13 6 14 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
C13 2 14 1.02547e-15
C12 3 14 4.03924e-15
C11 4 14 2.04976e-15
C10 5 14 1.20245e-14
C9 6 14 3.26631e-14
C8 7 14 1.66732e-14
C7 8 14 1.44119e-14
C6 9 14 6.83154e-16
C5 10 14 1.25759e-14
C4 11 14 1.53915e-14
C2 13 14 1.75274e-14
C1 14 14 4.10029e-15
.ends noa2ao222_x4

